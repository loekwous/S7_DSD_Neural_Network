��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�l�(���q�a��8`K�nz�w�V��� P�����"��l��p��2����}�iH��i�k��4'�����C�H-�%����c����ݮ�ƒ/L�o ��RD\���m#Ө���������tw��NA5b�7���ßS����2�+�X~듮K> �1p��M���%���|�8)�"���*q����E�x�-k��A��#����a 0�Ԗ~0Ghg�`,�i|v`����b���I���g �2|���KϦ�}U�+��t�qYBy"R�>D���tx܂�O3(�C�*U%f�[i��V�o���W�R�ѽ�	��Ǹ�L�8hG�]Ii��o�hk=t��zkC\V�P�0�{{M�^<	E�	��!G�I��E��/2T
�qd��HלgҚ������W�o/?Ґ���J|9�4��(:�zX	f���M_���j�)F���|�M+M+�D�j�eB=GF#�`FSF7�M��լ.|v��Ub��r[>?x��IOʕb�����5��X )�^k���q�����'̄�ThC|����Z�F)PjO�X�$4�G$sH~�u�c�p�������}y\V���Ծ!s�ċ��e7�p3)�c���H�V�,�+s����v��1$R�g���x��3	����tD���3E�[wI�P�t���5���#�8*`x�����=�m��e�)�B�gB�S\6��m��'<��#���bta2��[�9n gilZsk���8�S:SE��$P'j�������wM�X��]B�o[����j;^�&*�h��Hh��ł2=�#y����W�y�ʷ�Wd�7X�؋�KD�(gKJ�X�RS��{I��A�͏ЯoR���
�כa�p��G#nt{=���A	{b����m�p�^c=���Na�,�B��D��"��$��;���9y~4����nLܦT�G��'cُ6��8V�{������/3��x�۪"��/��
�j� 	d����lK��m�i��T�������9[K�|��GDf�&����ͻ�N�!A�:����_=���>����㠅��p���r)�{�Ogٌ�u���z/�ҫ�	�-[��TN欐"u�q[A,Y��
�dL����4r/�G�� 0�ګXk��o7����dXЁ����{�`��F��m
h��ܚ4{�C��.����P�y�wU٢w�����s�\��B�Y@w	� �<�񇅟�-3,��k����n
��I�4D<͍�?���:,�n�a�>h~���l>��<e�Y��b��"���g���)7�����@�_�}�:���+���z<J,t�D����Z�W�3K)eN͝O��!��E�|@O�n��"=�F�ɩGL�m�g��5)V2Y8G7�U&�:�i ,Bv|I��'�C��l|"՞KX��4�m�~x�o u��/d�����������r7�Iz�b�.���]X#%ԃ��QUeB�#�Q�-����o�O�W=�\K���`�$�ÙS��~Q�~�ǉ�0$=�p��6w�eB�4�?'��!�J9��iO����54��&4���?b�������RA�RZ6ف:�Л��t��v�����51-p�^EB�dkTF�U{�i�zޯ@XT�K�G�i�C�t4��|OKJ��B`ճNj��0����tPKZsr9s�f.;"��$)��Ĵ*!�Ust���)�g�3�(�%1J1/uZ�qN*�(@�M��E|&0�?vr@�w۶��H[�	�(��_>�t.?et�6��ߘ��c��j�Uup,��\*�?kBU7���$oUVLV�7���p�?z �Ma�JҔ�
�/�F$��Ԏ���{��V���#Y�⸹�I��4B2d/S�i�`�m�/嵐h¬���@)oXoVzV ��%�V��y3���X��a��J�w���t4����A)��DQ�����(XL�p>93a^������"kp 1oPbu������?X<b��YC��[	f�N�gt�
�BR�h$D�֑]�w���������k�5�K�B����^�!y�}����xس/90���Gz�/F�J�)��bX�%�b3?��O' ��鳎z���xF��1R��@�]@�	��e؄ݠ/��᝸�'x�J�fϴ����oJ��o��矴�Vܸ��d������ ���p���y�!/���E+�<|�h|ql@�d�-)��`Rrr��m�W���`��c3pKq�4{\�z��㋊j]��\P�@�kfъn�E�:a��JQ@��uyl@��X�Y^����rC�IE!u�(�y���l�^5�m4V�s�Tu�� !}�B״���t��)�J�oۋhN3��S�ax������廹�n�V��j���`i�bB�k�k���i�������A��_4N�$�B�-쮊F������9�qJs@����	?���JN�r�`L�����N��Հ�!UN�{�g�9\��#�߰� �PI-�ˈ�o��*�b��t<bKǚ��$QX���5��찆��<mp3S�܃U1�zQ��Z����t�k 0OX���,{˷g���j�H#b����}c%��G����o�%.��t�'�)9׍Kg��b��Ϡ:�tV�N$xK�N��iAd�
HQǰ�̋�<�W�Grb1��*tq���-�)$�u-��]������ 5ScE,����-T�=$�`j��b:J� ���I.�%���������:��j��
L-6�٭���^�a�^��!���̧6����@���c�3�4�~Ͷ[Y��WM�.O��GÑ����F`��Z���#���/_S�g�9�V���|Tt�o���I�"�	���E� �1��U	�Fa�D]�|ʉ��#|2q	�Ī0�; �b��4�y�Q7��Iژ��#2tb$dB^��I9�
�j� ��ĝ�QY:m8��;��Ȧ�Q"���?��~�S����m��F��K����,�x�t8zl�u��-oe�G��md���?uWNS����E��l��6�0��z1��>�প�A9�iޏ�e������CJ�������h�i�@;U��l��_�{͑s�r&gZ��dH)g�H>;zD��P�82?^ˮv�j�R>�����"6���|m'Tx�8�x�w�fA�Ut&L�ǡ��
���)[mT�L��6b��!L�<ZϿ\E��,rZ�O��Qޕ�%փw_���Ȩ\������E���K��<>��-S�n�xR"f�M���2D�k�.Wu���� Ȝ�.bj�3-݀Rua���]#����O��Ta�l9�����Q�p|���^TK�ͻ