��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w���N�?ƨGD$ܠ����!�jv%�ˎqʛ�������;��밇5��Sw�����;�7������5f\�q���U�5��5�y\��Q~�_C;�u����`��QA"�$1�^q˥L���F@̾
�q`�nf*�d�H�`O�,u�Re�;�U
ݼ �QX}9,�p�t���󽕌�#��_�NdOX�;V�q���v�����]��XwDˬ��8�?�͈��갱d|S�o,^Zt�f�CW���Թ�MC��qG�ǎ_�:���EM��/g�����x���g�f��7��Y��WI@��w� f�i��6������X�� �-3-�Ovb���0��}:�v#�>��_]U����1\ť����t]dJۓ���0u��ś�Op���m=�5���ٶB�t�m�	/�mW���J���m�cAL�\�n�z�S�H=~���mL�Q x�I�<�����u�¼��H���-*�՞{��MhB�d�"����|�>-��>=�"�h �+5&l��#�V�[n��J�~t�.�3
nۏ�SV�U&��ٻ�[]�C���Vq�j�W�+�٧��t�i@|�A�a���/�~��d$���sD�B�M���i�\�_Car�lk��W�8o-�K��$��_qq��UU�Ndݰl���Kƻ�!��Q'��~XW������Lj���b�gE��a^=K*V�3��Q�(�im��s�[� |�zC�Bg> �����4u�h�њ�����ՏgtW���T0 56��-n1���Q/�]b�
@^�4�K1���v �Vr9ޱ������84J�;�0%�>�%�cqNU�u���]��'��Z�����q<��/���K��i�C�UB6�MϷ�cz5�y��D�����q�/yI���͡�7��U;�����G�8dS�J&�\���aO�>��R$�����E�xq⟁	�6&��'�o�<g���o��q,�|��J��J�/��{	L��(N��ꊲ�'�fW�M�/���N��/��|�`���{eI���HßP�0��HW�f/͑J)o*+W!��~�bWI�!ӺI�U��������^ky?�G��'��v"�����p��>)��=�h��@�N��c�<	f©���4}����?5�O���^�A����~��Jb�=-Uh=�)4Ý��K���}ȁr�q�c�Ј�����y�	p-Œ@�]UQu���<~�t(k��	Vg����i����c�`5��~jW���1���OH���84p�o-rH�3$�o�"��ف�˹eE�{X��I邌� ��<��W������c{�k�X��ei�NVw��a`~�Q'^�Q	���
'l+Ѹl � @�_��,x���ܩM��m���]G��y`baCS~�Ь�V�G�����<�N��ߗ��n�h�뀨�� ��F{���V�%�q�Ӛ��Z!�2�D���Di��%V'q��H_��G�_��H�`��������\,�[4�"��b��� ��^B��g��Va�Ez�_oCn�ò7xc*����󱪓���W��|x��魃�R��W�"_4��3"�@j�Z�&Bp�@��ڶ��_�rM�󰋡��E�Vic<1�!̓�a�Tw@�)���1n��{��:y�#h#�c�JT�'a���yU��<��%��á�X��7�N~�<��t��c��Ä��R�q>�L��]=�,�}�+�/Y��o*�S��e.���+l�f����}� C�$�������X���5"��
U�� ��hӁ,��2 d�XP�Vg�Eg".����0LW���mBII�MԸB�z·ق�G�Y��ͣ>Wk���~@�/M�b>�-2ֆ�ؙ/2��ŏvo�P����ͶZ�����j���r}����^��������=����������W^��B�koEU�4Pi�&�� �[��4���u�8w�e類X-Ĩ�ZFUv��әXȜ橻,���۷vnB9Gf�͹EXdu- I�+��`��\c7�ڀ�߇taN6�ȩGa�yDP�'Xĩ+��[DG'��_�D�U��Y&� ���4H��,����$�z/z麑41��ڠ�t�	^�[���NQ����a���S�~��|���FLP���R�|_L�y{h�����JPwk�=�>�� #��C�+�yDe�!��׍Z��i�N�cݪ��l���>"�,1����:���~kh���痢""�b� �wb8�7u���i�[zIp�/���϶�u(��U�߆����.�)U�$B� L�Zg`����<��^���rBکЬ��q��z�����B�N	�b@۞U2I$[��<��`���l��u��g3��t��SP���) Y&�ݧ��(�{����8xuk���D[�+�Q�$O潰џ��	�Ҩ���n����8�L�h���.���+2CX�v���ta��C�oV��"­�/^�"/dF��G2@��:6���-�Y�4$H{Aè؈�ŭb�{��n��րem��i�]��F}u����U��J�6E������%�B*@� ����������᙮���@�Y��[Ax�PPCI.��T��ΐoi �������"p���wJ1}���,�����ǔ�LlQ��!�aߊK5~�^?`����j�n-���z���0FǇ��iK�<���"b�+8$h�����l���k̹�[����F�LGi�7�e�]<��ax�T�'�YV�0����9qb櫃x'�{�v,c'Y (<�����J*��������S�ɝq4ހ���2�.s�Ih������J���"���s�w�@"�.�n�KMDr���J�j��=W[��cY������������3�[��]C�o�h8<c\��Ar\�ԘtK>,�b[�q N�5�wj�=�r4|8�8$9��1<��}a��Ϳ���}pqQǗ�X���M��T :�B��*�E�(}ɏ,6�?ʝ��q��/;��f*��e['Ԇ������_��c���`�X~>��o�2���y��W������˼@�;�~��:��0[U��@�aT����BN�|�6h���q���ݟ��m�6kI�x��77Y�����ax�I���-1�Vpz��D�,l 7锉lj��,�y�xҳ�$�hŞ�[�K�w~�bSVv0��&�;���Ʉ	�t%o���Ӈ�=)��s��(�u��|g��r=��&%�^򄖓ֻ��h�����H������Yt�h��0�=Gר�|W�	�s������cW?�i̹d�_����E�q(�}Xk��r��VV�Z��OK�:���=2��[XQ�	4l��;>�Bcd�y4�ƌj��	�6A}�RQQ�L�H���I+����i�h�@Ai������K�O��J(��f�{U��o=�4�����mjR9��P�5ҧY�c�S%ı�à��bA%L'Q�& z�Ds!\�,s�"�9S���Ǘ�Z�� �`,��Z7���"~�hII���G��Q<+�ǎ3o�bG�zb�٩TLC�$���bV���G6+� ͇�f��w�pL�=���.���� 4��������$q#�Mf�C��8���r�(u�C/�~���.�)&� �Ǡ���� ޹��>�$�6N����U�-,(v9�"�q�i��RO�
-��X���V2�(֚�������h੢��t0m=����0X;��R
 >0Q����{����2^�Rɐ���H�e[�N�͡]$�J��mH����1Z�(������]���;Š�ښ_^>�+R���?ٚ
&�'�,�<��Y3�1��E��,�b��f��� �Q�g�ZDS��Dʬ�X�&���`B�h[�V�^�����V�[1��px.�*�"������e����_���բ��q����BL��i��*�ŭ�=y�Ea% ��*=b��8�*�+q�ܤ�T2w���C� w^���]PP�$>ƹ$��|͗<�ֹaG=�b�O�ͳ��O��r�g�y��.B#{y��TD��<QTsċK���s��H��}I9�$_ ��d�dh۽��)7��͹��l9�3��uĶ�ډ���
��d��f��#,���-r\�?ّ��U[;֚�1)�w�AY�E�/�Nذ�xӱd�{��܏��mP@��:ǯR@o�Ox��3�c��XK��P4@t�QJ���䋒�_�Xǥ�ªU�0�߂��-䳟�\]@�l��X�"�X��)�N�b� Q�����!2g~���
~/Ku*��ل���"]�����!1��7zK�E�]Uʩ>e����ʹ����+��
:p#{���'�Zt�@�Ϥ۹;�$�[Q��6�f�5u/u���{@��9�t�)/�l��t�3,�^@ˤ�M�̈�_���q��]�tx��n�?3����\����WF�x�뢔��h���u�0�ρӍ��i��y�N�:��
���� 	Pb{\F�˿¬��	8��&6�K�5R���<M芄%2��Y�pCm��5ۮ�=��o`.�7"��Yۇ�Hb��4d�O��O�W��.�B�U�yk��|ƆhQSa-Fm�D����_��7^G6�d�Rwk��F܌����no��V�JܘPE���Z�+��8��0�ĞѦ��Q�����T� Ӻ`WO4��6oӨ4��x���j���|��?��<����rI�B��G*��da�;��(d�
��p*'ߐoQ��u�;�;v�LZ�vJ3���".q84Ґ>�����;��e<K;�g%$�T~���Q'��6����2��j��E��E�^� 0�@�����RNqR�����q��Ƙ<�ܳ����"hm���
3�d��[(z�����¼:���
�і����lيaSF�q<��/�8�o?� j�_�|�ŝV�ܼ������yRc�w�ڦ����]�=혈�Zha��I��>���~�WACt*���D&~�?eD��@����b��>K������F������q�ǌ����{.v{C����-{�F ���6m7i����E��os��ݘ�ܭ(�V$�g�$_�v�)[b�v�����-��HT�IYWм]|S-E��z�q��gD�N�.�:��� Pw&�]r��/�+$�e#��M�R�K�W-�t��oZ�s��~��)eW�E>���#'Ѐ�j�/���)�s���v�I~�{�56�Y껨�z�S\��Nֲ��[�"��W%��<�]�����w �\e3����ɻ���SZ4?ZdͰ��4Q�f1��(���+�	z3��SC^�{o���}4�m.�m��=���҆y7�J���Ս�D�:��F������e��W��;��@�{��VQ�Q<�b쀆�p�1X%�v��.��Y	�����	c��?��I恆����K�.���mB�k���J���@�nd����	o�Ȏc���Q�]5o�%��s���][��hY�|��۝
w��:�����qH:2F�;i��jw]xm�!���TwF�co�&�Q�χ1Lo�ˈ��9B�Y�\��?��v�e�4V�u��<p����z���U��m�@S���I�4*��׌�����51��1�:qb�V��LO�j�t���N��[��V�\>%�8/��q�o"�UI��[[u�ߖt��-�J����M�iA'�p[o�ډ����$n2+k�?� ��;� ��/Qe�G��s+�`�u����٠<��wLD<��]�	��T$�*%�N46�����J����ɷ
bGjAֻ�\�~fUU�l0_��I�'�+8&p��@�5���U�I��/�9��vǥp��:�#͂�ƃT��*���G8#������*^�V�U��{JCq�������G���M����qLmsJ�h�#����ۄ?��b���O� o4�
�� B�+vy���kc�Q1�TW�ug3뷒�����a�,�>���ǤTv�@���[�N7AfL&YmDx񗒜W��h4�V�����*��|��G{{��8���ܷ���Um`�B�!z'�sG�a�xb���5��[���ŦQ�q9��m�&\���Q�7Eg1��$7�5���##����� �B��
��)��W)dA�'�r����Ǉ���g����&�>9~�7N0zר8Feg�F�=�b�[���CS��o}j�[9���@ȕ����Wǐ���FM��lE���Z æ�����W����?)��g��u-Cя͂2ˡҖ��g�1��>?��M��������T^�w��<4�Q7F���ӿ�>�g;e���'e�N�����9ڝN�C�ن����ȃ�
ǧS��f�+�$�`������g�@��p�/�'l���Ƶ��S ��i��`�!�'�=%��
��q2�-@��L�������ZڀB�Vnm���ݝO���]��歮���x���W�b����)��F�J�ռ�t����St��"<�
�[�M�2����j��ʮ����'�߇M�U�W"��0Y��~�v= ���t�?%�ϻT��#���> ��7�17P��� ��������-_z7P�P�g��M��i��&�Q��p�����(�XǍ[>ˊB~��Ĝ�]&�5�tQ�d
X�V�-����A�}v���9�`�#��qs�"M�.p���ݪ�w�܆Y�5�С�2���s�L���G�b����;�<:y.zE��aP����`��m"dz���c;K���>��	�*�cA�y%���a�hH'�L���s��q���N�*��,�Ϋu�8"��S��q���F�/��7��b�8UQ�%��u��+suDLY���}ޫ�h�FE����L�3�a+6L�i�m�z�c�8�T}5F���n�p�����-���Cg��	�CMn�Q�@YQkr�߬;�4U��.��Aҽ����8�߄��Pߚ0+�M�`�d/���Ӎ��ZQ�[�&
$k�3�ڥ�<��	��m~a��y�]g�-o�yR���X�*A �K@�t˱`� F9^����9�1V��ĕ��[1�*Yϐ�P	��.�ậ��i@EU�M*�`#!���ɳ�«h�HJ���V㺛�Y��ڨ�i�ϜM�����k!��;<$?�IS�1�YܓO�`a���?i�hqs2t���o��`�J�
��&WG�����nf@��m8F�N��k%�q:�m��/�է��C��|g����9���]h��c����1U �����ۭ��F����=I,�ۼ+��lxNM�EE��f%ꌠ#�Oo��ҵ\�7�5��?�k�]ΗT�þM����.41z��/=ھ�.��󥸘l�M�q����l��c����ءB�,�鼯D�<+����wv(4�F���x�||ir�O��?k�G�͕�|B��L����u��������n��T�7CPJh�t�{{p�m;ULwis;�$1�*��=��s0���w`��gKl�5��}sb�]��7 �#��G
j]��N����HN>�60�
w��<aD ������_H~��;����D���R�A�`�O���M�kX]��[GHwS(an#�z{�����t�Q���C����XH�\#�����~}B��ae��}�[�|�>h1*R[�}�O�(;�#������ܴT+n1Q�7��JH�סi��Ȍ�����@=^�6�I�ߙ��&A��՟\�^�
8GdJ�3'��%>9F'* �6@�t}�����߇sA���*�_ *���3U܊p!`��>@4k86;��C�./<P&j<D70pe\���D�N�%��'g�d�}��2���k�u��L������\������8#�%}��ɓ���k�Od���`@�s.��8;�7�*"�ю��8~2�N̈́��,o��4q�EZR����k���Y%��k
h�3�T�AUP�6�R�.[cR��u�/�+��W�HE�'�����W)F���0"�j��������t�QW��3�Q\�٪�1���U�!��xͶ��pM/砽W�m�Y��R��K���bt�O���Nޗ^���ʷ��Y�UP���Ī�����1H� � �{ 0�X�KF9�N�j�P�i�����Ϛ�ȃ]��/�W���%TyQ�ș�²^g��s ��a6������xA�����D�ѕI$v����pM���]��=̷�GO�:L7Ld�R�Pv��9��yO4m_p+N��-����|�����z��ׇ����m\fO0��t�6p�Q�5�WDA�=��;3Q@I�@��=