��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��ӡ;h�>�C�0��̚EvW�66�Q�������:;Ra�z>#	�ɶ3�=r�\��@�Dw%ٕm�pQc-Gm2=V$gP�q�:7y�z:{z^��^Ux��wZ��#�Y)� 2�X�q�+Ş���dA*Q��(#+�^��w�E77�?���/�V�t��k!dM43U �!t����h��>u�N�/�#�B���*	��~I����]�s8�N���3��\�GS�����Ry��S1�{%�V��k�ʐ�Z�L��ȁ"Z\
�����
�9N�b�/.�I�в��9I8gm�Vj�����uB����B��Q���6!j\���8��ZV�Î�f��Z��Z�mg �����K���N4�Їuj�,�S��m�{��{' \M�{Ú
`�����U�̓hi�i9���ҷ��I��fB��+ųձd�����]%�ay+��I�癒�exU5�|��*�Ω�^d�mb�H���XP�1��?�g�dU�t�RX�<aVa��J^���� $8Ι���Z\���s��VU��:_�{�X�	�u����b_�r�!ia'����?�� �ILsܒ3�>�Vh̿(��*�?УOT�eQQ��Ң���՜"�)��q����3�O�S��%�th����*X�8�,��-�=%��ɂ)� Y�%P�%����[4�
ؐ&�E�~��n�}j�o N�]��a蠾E�I=?���5FOY>qZ#�X���'�e�o�/8�)����4%g��I�;yO6y<{`̀�*�Ӷ�!��\d�{b��Bs����8�\b4����^�ńz$Xζ=�5��:Zl�=?ĺ2[���r�R��-1i������N�ou /dy�(�Ldy�?��D�?���7�4�"�^^$�Y�E�����X��u�e��Fm����x>�������`ڢ5��^w!h���D��K�g��.��~fU��6�R���{��"��ӟ�2��f��|P�����D����E�7P0�	�t^xɊ$V��*l��H�MZI47�>ĕ��犒%/�O4�d�W��cGq��}�(\�qJ�{�Ã
K��K	����9�>���ˢ�N�3�%�JPY�uJ'�ݛ��� �]|u>m�74J:���J�:q��c<����V���a�1�H�)��2�(0�ðx&^�D���frA?I���	�>s����r��c��ͭI�]�Q�u�A^,��#��)Vk�|�sW �=�P�K>i�kO"1�}?���8ըr��m������V��69=i�L�SG�����Ԥ�!~��R���#�R���>O�q�����!�1D@Y!������i���{+�#��M���g�?����[�D���6|Y��k��4�*���a�~�-���#f����?S8���--��U�1Pwc%�Rr��է�f���
��f��Yml�P{�]^����<j2fv|l�Q��u}��Xp��K`D~�L�d���%^��L]��iia�X��)��n��#9O��d����l�#��V	6�b�V��CݰsTł�#{��>��ôP�N��u������A���`�,�(QC��S�ϕ��x�>P$���S(,%DC��*l��jػN�bӞ bL*��X�t�F���vEh�a�~��/�X%Y���}�ќB.��D'a/T�}�9Q�(�jc���DR��"�>��1S<(ۚ���<u�֍Ӕ'��_0���ܾW���O�6�Jf.-J�q��=f�Z���(K��@��
7b�����ˋ[[�ʉ�~�E0Lw�\-�kf�Kz��mR�n,�e�����R�8<�s�]�������@�}�"����=�8�&��r�E�D��|���\�E%L�X��=�_��K9�G�i�rN{�(��,�<Й'�.�|ko����M�j2�_�UsfӃ��� ��7�i�{��?�3@�����k�0c`߹v�$I�Ӡ�Uٟ�G%��*�?��!�N��9�P�\{���s�ށa�����>��=�h�Qw
�ݧ����C?w �F�r����'�koȜ�l]N�o�k�� �c��Ծ$,L�5�C8����.Bu�e@
@@�;6���wz���A{���E^I������J��!_	P�B�t~�Uġ"��B��I\u�Q;�f��Ah-�<�&�-@��e&�v��id�o8�
��c�⒠��1�m��c����Hm����e���96�����M? X�u����e{�%}[�4���@�D_�_��;�w��*n�Jfr;��Q����U.'�0��h�i9��QSV	Y���XD{��\�z���u�nld{a_��C�b;��gO������'ot�yFHҀ���{,[�W5�\15��6�OI]�Ž���-ĩ�!tĉqgڥ�����}�އ`e��]��%�J6�����b]����K�ڋQF��}�*4*��g�D M>h���0� ~�*� w?&��)�)k�#g���M2��n�Rԓ�����ma�Ԫ�(�0�,?d2Z\�� d�\��P��o���D4���!�4g�n}�j������u�IO7�(W�C����<嶱Z.�Jq�|rA����Y(7�������CV)>���ě�lgRE�����i�g,M��!�4q�ݓ�Q��u�t�RLU�J�|�ą�B�&�uq��%���9����������rL`V�IuA�b�z;p�>�_�1��8���e�Eߙ#����M�������L)��������[f��xA�4}��V�.� ~]�a�2�p�sP]0ģ9؈�U8zg�E��X�s�{�p/��׋����<L���������R~�N	�	�·P���A��RP
�$�o�?�R.N�|q�KU�+:7�������ӟ@����������%��cx?�:��\���[!����k/�������X<���B|���OT�A_�n������v��r�ȏ_�ɞ;hN{��-�����S�U��C�bk��T�j�ZҺw��L::A�5�������l��\��$c��߉�R�E��EP��3)f� =�SeǮs~.#��|_e��������T���O�\N��ـ��~yh̷ʤ#9$ڳS��O��E#P��ȍi�)Q���� �V�;o��1ŝ^�ë�ڽ�C#���2O������0d�g�1�f�ɔ@���c[��u�����o��K��\�4}���]��lt<���*Ҕ����) �J%�H��MӨ=��j�@�R|�zN����~�)'�����`�g��dVRA&���J=��M����b�`�
��ymz`�9=���_�L^ݽXy4�}�CU�uީ�/R;;�;K�{ ~e�V��j�"h�f��g�2���Z��ۂ]J��;Kx�)*x�h�`�Ojq˛2k�myP���#�� ���ȉ�P�����u]�3t���to�-��̒�K�Z�	&+�Uǌ���:������ ��ى|��ƑX,{ŶUS��Ӈ�����t3SNR�SR��\��+�5��������d4���-�uPzZ�
;6�|V`h��G^%���TV�{�\5˷�ȝ���V(�;��������>e��ݹz*;��#�u��j������ސ�/F���A�s��@�4�� Р�r�l΢��G���%�$N<���w��i(׭���;�%+ջ���m�9�q�SI%)��4�mż���N���V��JǊ�HTד@:T��8�BOځb+M8�^	i;|�Y�D	�P�r:���Ì�>ED74��8��-�r.:�#R-�M�"�o/d�o���豈�"#Q��䫈h{��?#�U�o�nG�Sj��ǁe���Y�[�l�B�J�e�p�=?�eQ�cr��	*5�g�Ju���	)T�cS��|fFZ|�]�G�̯�F��B��|a��28��Ӆ\�*�x^䨛d��;���[�����3��b Fl�P�S��}-�z<�  s��6��_~�2�E�';&�ߏ�4����
��|��^�TV�i)uj��s��>�p�/�t��)��.��S��n�|�6��gH�f��H���J�M/���j�Z�z�������㨞Ky�1�G�k�)՚Y|�tsAV�%%�D �;�q`����U�������;t��� k|��+2��V%٭��CL0{��X�r���Y�ܤ��`'c(.QCN� ��o���Rϟ�7���d�t�&E`Ê����Qwc,�=��3����Wʫ��f�{lp�S�+wޚV�O�}����Îh{���b�X��ke�u=�d��9S	 �|9]A�3"-����</��#�K]>����p�� Rw,!T�܍�t�Čk��uN���F�q�u�E�4�C� F�hGs��?�!yw�۳P�rb��esW;�m�;�	�-�r=nLd���A�t��L�����aS4�R:-��N%�)e4U���A���1�v���9,�]��<����B��*�q�</x��"ި-�M�� �&05�_�Wҷ�h1�p��l�{�0<�4J��_E}1Mx�q��ڲ/�ȴ�4)�H�m�p��p�h1�"��:�<�J��߄�C8o�ᤃ�H�֠d<3�M�8��Z��3�@��9�]T�9�3�$�BO+��a���'���%�  ��S�la�[�����g3�P��j�w~�yk�^�7���*��v��~Ό�I"�.y��]���t���\�V��a>��%9 mr�>��{>�[7��Y��b6�k���J/32L�4Q��.w�뱸�?d�qU>\��؝�}j��]�$�����?�Q��択�����x��'��ͧ��3��M��(�l�1~��x�a�����ᐾ,����R{��e ��3a`�/v-�1�o�R�X9��\��X�EG��U�mA��X�{�i#�S��;�[�
Ee�a�p���)��k�
��R�b8���k��j,�=�@l}.��8Qm���[^�{��'I�v���L)�fB$<ع���,�\����T���QГ4W�V�N@2�V˨R�4�Ů�Ԍ�kI⚳�����#�-Yjk28��Y�5E�7*�c���S���i��g���R�I�A������ż�`[�Uܟ�Ha]�Bkj9�L"���3ӹ_l�S��e/J���,�7/����bҍ����zU��'��HD�����J�9SJ��h}m�P'�z�!G{O�ק&��3�� [�J{��c���Ca����3�lf��-�;�?�jWIO�Q��7ޓf�m湞�D�Qz&l��*^�Cs�JB����.f��.]uI��\�jX P��`	�C����?��@��aLK��'|��_]�bC?�Q�NN�n3I�-���1�� 4���}�QbPr�G�O2������i���WB�����/*L6(�	��[-�w]�#�z3X��E�Xp��Ii�v +�n���f	:�t��D��Y���
G˃�z�cy�@}�$�ACs�:���v��J��1�����c�_nꓓ�u*{�{>�`nW�N��T~�$���'���Y�~�dt�܁ ���5|�PHkۘ����f��c���������>��%���4S�T�i$t-᷐1ꋉ��&n3�bx���,�7kH }�Zg/t`��ʨ]4����� ���I�?0{>K�`0�Lp�xF5e�2t�|�lfڲN����(�� ,�n�Q�h�=d���5��Q��tA|�@Ub�R�^�@/��X4���,D<ƞ�7l���}����Kf5
7��#*�N���ʇ��|�<8���L-s-��"�f�!)�ZM�rs9z�hJ�d^�ڝ�U��"M
��e�>ҭ:�+Т��8�kg�U:lHED��18G�а������	Ѭ�r���(J[�H���T
D�DN��s�]CqY_�y�bnh�[�@��7`%�R4��U��4�!�m�3�͟g�e\K)����d���p�选Q[;ro���1��yZ����0_�^�|l��N�#Q5ɴ!�����n�4ް?�!������X(��I	h�C�����\��$�z��Ka=Ǎ�M8���@+�u���^����u#j=M㉠����´�b�x=g�����W��n��� �U1ө�LB�	��i1� ��+ԟ���݅�"^����g���P%�]���2���i�R��Ps��&�/�>fp>��gct�Z�F�~ѦO{�UV��( ŭ9l����
���6ŕA@TDL*�g������\��/I�5L��1QإJ�/Y���"XO�p!�ZE�\裰{���3!�Zm{���k�+ϺS���r�1��η�����Gα���w,V1��,/��g���d�a�I軾��	�5�_##왍��C���1�H�jL�a!��0\�0^A�I�)|8=�����<T����mG ������=��Xo����*:Z!��g�����I�"5Ecl�����@˷h�`�QgJ0?�?XX������x́�3���x������,����_s�+���ן�n8mjg*�d	��U�5�?��p|S��b!)���CI%�)�лE�iɋ��K����gk��;��L'0{��!Q��c�|��ܱ��㞉J�>��[��Ԁ��ko��[��:� b��v6:��1MF*�:��5ͪ���^wK�(]�A��[��4��B�BrmZ_������8�0̣�G�#w���k*H
�5���?�T�s�7V���|�V��p���"��.�ƆG*���|<���}��Q!�ӃdAu%�[��Q�~;�\xݔB�+2����o_߳P�	�r&�=���)�@�K��$�46f���,c���*G�k_��
�j��-O��a�/�&�cu%�G�,P6W*����X���^f�p������q�H�bwn7�T-J���
�>E+��h�ew��"����t��f-��xs��/}{��w!��h�87�!�1p�-~�CW�g��)�Ja�{ßSe�:��J���;F��.Zwl�̹�PW��u�OFW32����8�o���l�v^����m�u��T�dK!^	 U1w��B	���U|"Lx���Oa����}0^A��K#�`�����@Ps3�W�$�d�EЅ�U{�\yV�=��$���"�NF�6w����.I�u�rw����%� J+	���XAӨ�MWa�q�Q��}��X�{aDi���MP1Z�~8����;h��rE#MnmYP���o_����\��׸� C_J���R�F1�>�dS@�욲.���{��&�c�6c@�������Q�x���#�ų��� �x��c���,!�@�����ḇ���腂��v��7��N�D�J�id�	HP酅�y��!�e����R{T=�b\ �bKb�!w�l)N�X����F�������]�:F�7{\2�Q���`ƶ�"�yv�c��X��E|�u����k*k�
ж^wfB��3�:�+�z�Ls}p{��*���C	hV9SZ�$�t�}��g���;���zX�Ik(q�}���e\V�JZQ��8�/�Iϗ}"��퓣�^��&`�y��j���^�f�e��&?�����f�ߞ��%#�A���)١�4c�T��E�1����$����7�gn,A���rR�%�j�څ�8�8�[��uS�\����FU(:�~�H�}_�L�yBs��=y�#$iS%�@����c�?{�¨	�o1�Rl����k59����3](AȿTƾ����#mD��C(N+��9��a
-���|U��W���sVK��]���PZ��sF���?�[�|������(����b��vO(�~6l�LG��SEi�Dk��,#�Q!����%uOI�e5+�z�w�-��8)��.Z�P��.�bt@�144���4m M��#\;�P��}��_��o�+���1�A��M}�$O�Rg�䵻G���m�d%�xv/wm.aڳ^��z ������ ���*g�>wQ`ˮ )�5_�aI����̺޼`�g��W6�WV�n^J�{LN�>�A��^���S7k:������oم�m�����hCB/YY9�F��	>/m#r�R�HP�C�/�� 4�'[6�"�A� ��pp63�M��,�2��EݯB���p��H��P�(E�؎�}\j�sg8�;�_� UT>�#ʁ���J��z/X.�I](�';�-4/�ly����r�_���ܸP�p�5J��vUFN���Tjn�˗z8�v+�f ��?ܿ!qQ0F��} ���yϛu8�=J�XO||5��7td�EOe�����GxJ����H�f�6m[����N=]�7ш!�D�8����$E?(��8��3�Q����O����![$�Rp��h\5�=)��k�E��!�(y&y(�;V�U��I��3����h@a�1����  R�.����N���5w�Ò�u�N���[���G�$��"l��SnA�R�����s{���4|w+��*�Ϫ�s�,L�w�����(�lyn!�p���1)�P�M�)R�5�*{��q��<y��&����e֕�qQ���k���A�`#�o���u´�@���c��Mت�ِ�?�bd��%��oZ^g[T�kdZ����m�|��^1IBz2��^@��pUZ"�����2����1����)�I}&�
������ ���d�/��4�-�Gf��{W��y�I4	&��g���3�<w��4��D�����@X�z��dC��݁c�(�T����ǒ��;vR�F�o��G��H����LI��3%��̕��1����d�������q��CЂ�̊�?{kNF���f�+�C��Tm��P
ފ�yB%2:M����S�rA-Vv����(ׂ�(mfGI�d_��*�����9�4'���9�g�׵����>⾖/��-_���dѻ@�U>xuJH�):E/{�DZys�]-ċ���>b}Dz�h��JW���u�<��<%��a�
~���|�Uk��X��H��Օ
�r��3���Ym��S9�!� 8z�A��2�|gA���4�����	�+�45.���gf��Z�کJ��ْ�,Bx����J!P���-�;:�1�3�l�N��U���<	��-������O��z�7J(��b�z�$lŋ���E��@��~�ײ��t���Q�9��-^�El(�}Vt�R�W���jh�,�ZO�^����oxif���h٦m��5 cC�y� dWA�Pg# j�+������	���nC�ӂ옦\��z�rG��$U�L5`�7�y4P���I��Ҝ�y��aç&§l�u����c���zK�!�������#̇(�N/Ɯ��I;xLJ״�t�5k*@����­�'��?m_�(���_Y0�p)ѺW'
�H�.i2h|�_nv�p��I
N�"M��f�^��W�Hڞ^�-�qD}�1җk�p=�N45߁[$:z[6�w�N�q}J�䮊�	z5�6���%<��vW+ϋ�o���d ����Qd1� ��LL�!|���M�&{<Y��Ds&��.ޭg(��3�@%4��s��N�ζ�`��Տ�����?!�h�k(���$��A0�I�z`�^���%8_�������Zi��C��n��t�)�c�=�󮭽������y�*a��}�ll���q9m���}C�L�|8�#<Y�Ja�j�g��@g���b�R�i�PA��;���/�]�q�3�K��9b)�E�#1��\�C#��+:/&�y{�u��U�	Vg�4Hp1�<h<rng��Q��z�h�
�=~רR3a�D4� ��zB�����oZ<+��s�+�0���F'ƚ_���c^	�ńk��H�,�d+�)��Z b�=mx�''�gȕ�U���V56Aĩw�����jP���!:�����N,��ԝ�U��K�%NI�x�B>�A"L���kV���#Jԓ���[�v��Y�\Tn�f��+4��{���wKv����`�Nr�+kը*9���[��=��[�O�����B��)������n��S{��6�X��֚��e�ǉӜ�<�W�3��DO�͎�ǎ��-�ܧ��c�F/�j@�\<	5�k����p&�Xp	�r�ӟaY����ڢJ�Vb�!h��<b�8�>�hj��@ݼ=�yX�@�SPi���`�p������e�6%���X�d�k���c�3
�H�/�;u�cl�H��`�nI4*b��7}���k�r�O ,A��_��X�*/œT���	�I�w� q�nF4��[��B2���6���?���of3lR�Dou���8	^���V0:[�V8�+�ߗ-&�Y�I;.���+Y3q�JLi����&�[��2����,�!7���+P�:�F��Sߝװ-���2��g"z�K��B���g��,�o��bڣ%�^�3
�+-�b���C���	1�dH3�$f~YkjF	�/�\��xA!"�k]s��_��P�����*׬��.L|�]�|�����%b���/[ـ3�0B&6�%#{����:y�:*VȚ�g�r�� ��D������!�
�d���o�bG��8�q�������&sa~��IF�F�6w��[/�p7 �|���Y���p��H�֣���%97;�t8�)lz�4o��;�߱,��\\%<Ʌ4q���+T�p�8��o}��S%�4��̢������Q�u�)�Xu��A>�^ȴw�Ft˲]:A$N8�d6�jbL�"o�`�ɒ/Ë�߰QmS-�_��ئ����ٺC�:��+�?�ÖZ�Y��:����LZ�=sԕ���#��I	_[1aB�L�gJcAM�K�C/�(�%����aS��~YO���nz�l�t�S S�������qE�I\j�t,�=���3/��Pѹkc��]2R)_1V.�-#��2���MNt���Q̞�M���������R���uX��T
�ã��WՒ��������^F�5���@_e�������0����_�s�x�Zo�^��>]�e�T�ڠCa:>�Qy�O���ο��Qm���@�A>3����'��"��-p�&@�6e�X��	�_*K7mw��Mn���_MޏN�gClQ�ؼ�H�*J��r-^��=du?�����	��2m:e�Y���%=@VJ��I��J��]Q�ޒ�D��)�&e.�l̵���� tU���u�+`G9�n�o�7��·㒉7*�I�/��[h
)��.�`�8e��t���UΔ7%�����ݺ	Hā����sIY|W����y$w8&ܞ1q�)�|�F+�:P��Y;i]0��F�/�ɮ�߻��πM��,��B���nh΁L���P�b��J��\�F�l���*�K&Qp�v��9�N�O<��j`8 +�z
�h�n�H���-ڛ����D/���6�ߍ��7C&8���AA��QtO�0�n��]�B�C���O�фs%6;��{�Sp�a9��4��A�8��v�E�)�-2��ͅ��tck%߶�;Ҁ	ZML:��>�.@FfF�C��� �梇��Lp�?��V�@RV��^]���K�Xj�574�g�O�7����d��?�B�� G��e6�q��}������\)ӄ~��~;m�<��2��0��m��\g�]�OLK�>:}><�������{������k�g*����b7y�3E���R1���0ʔLr��W���5�a�ſ��4?l]�<^+�<e�4�Y��.C��k����tB�る�.�7*�G�I՛x��Xa�77Sg3��X2Л{+��ob-Tko>��Yx#-_#(�~Տ���/�8�!�{3�a�m!�޺�	,�u`��*�����OJ�z�
D~C�HR�G&��u_�r�N:��\���?԰dմ<�5^9���5���Q�w�Xӏ�ԝc�΁kR�;�W:�A(����`�W�1��ᕚ	�vT��uY7^FT�-�[gBl�2�=+CT�P=nM�N�#�m�@�>"�x=��6�ċu�/ȡ�r�;V2�p�X5��
�� Cx	��0��"���Xh��Vػ���H��	������Jկ]���'0��2�A88�r�P.�yט]�Ӑp]����wr��>�S�?�l.7 �)����*��F0j��c��L���X�K!~4h�?[Y�̠�x1iy���%���O���Þo�'Y!�"D��f���f�/�����3�I�>���/_�� �`�����YF@.���Ŕ1o�)����A��i�@;���
D��O# ��7���#~��!L�~v涥��l*��U;:�,(�&�C�R�V�<��F���h��E�d	�m4��JC�FZ�aF!d��7�`��i�O��p���ě:�A3�&�Ӳ�*�����MX��d���]τu8[Z���mX�H���{p4Y�� �CmO��;��Lm*�<�!J�$.�j�A�#u��t��Y�Š�"��<*��s�}su�A��d��w��H��%�{`����Z
�v`x�����4�}9�e�꣧�FC5G�f�Y;b�5%>v����κ8�
����j��3�Y�DfMԧ)�1���y3�Xo0�P�5��t� N����.�Ih��?9�Rd�겎⠠���3Ǟ�%�b��k��]=�����u.��g�������i��-��)
�	h��R��HZ�1Uը7v�G�2���[y�#.�}S��Pz�4E��(MtN���!�����GE��b��8��ߩ7�IL��c;����Ͼ�2��3n���o�l�jez���9�S~�z�bb3�*:��E3��-=�WV�@Q�l�iH�V�CI�}�|�,����ݔ��CƦ_Ζt���JS��Ҏԥ�w䙒JF7�����cc�7κ+2|#�R�t-� ��r=���������<o�� ��4c�������؁�� P�>�~�V\)U�U��;$��u�`oR1)�m�VqD��1�Qm�������zi;.�C;������8_�&v�hpos?*��#����j�g
}s(u��'�\��2��-�B^��0 ��İU4�i�4�9R�4��:UĴ����Fl��8��yDG4FBȖ}�K�Tq6T9�9hS]u5��G	�`�M'�N�O�2�[+�R��B�P�$hi��$��%L�@{l�Y%e�l�h����x�w�E����&�H�p3�o�-��Q�$ޔ>Dn��u�Br}*��h��,������8�����	%\�X��S!�������OlPh���� sߡ�|ѐ��*�+2�Әs�:+N��&��n��*A�yo�ث�2��a6�p.h3��ҏ2��I��͠��P�/��܂>
�D�q�K��ҕ,�e��i���s~p�[�{>�MM�D]J<�.��?��56�u�5��F(�>��2cb��[:xݏY�K؀��I��tRY�D��&��M�tZ���ӉWeq|Õ��.���e��e���A�@E�J{�]���)rNU&'@]��4�ӗ�A�{h���H5���� ao_��������������Gn�ݝ����a�}}|�#Ơ�ԑ��ưk,�˳�6�tmb�������l��:���,z[���,�������ꃴ�*��_̵
fҊ�
�������!NthC��Cq��h�������u���� 
�1�4L Q�����';E|��RC�$��A>���e����A4�h�� �:��0D=��;�e���6���դv~"\��;1nv��L�w����蕪�1������}�g�獿�B��Q`���TJh�:u����C�� �k��4Z�㐲�[�ɛe�M֨�Nx��Sʹ���5x�F�j�=B�9����x�{N+nP1�k"BB:9,䬞Ӆ`V�&��dB�z��%�r�OC[m0�|�^�'�ȴ"�v�[%�㻊��a�W���l!+���g���+��c��n��(
��L8*"������s$c��6�Ʉ^�fZ�H�i�=�v�0���5K��OB[�%�raK��;.�C��AM�����Pe����"Tt=��J�<�rQG�4��[�h�'w��|`̘S��e�+����/��cɖI3c0�WF�k!��V��հ���OmU$�K5HG�FN9G�Ǟ7���G��� ��e5�z��ݲm��!3$"m�Վ ��L�8�VP���Y0}�r�����1��$=OɎ��T(S�>�n�~k���S�jW0ڣ�x@;*9��Mt�":� 6'Ϯ��]Vg�̡�hX�ru.�%��)Byہ��f�5<�4���R5'��;g2�?�ۨR��~�����v��]��{5��eמ��;K�v�7�	�?�Tu'���b7��P^l�[�K��"K��&{�9����F�4k j�Y�L�FY�|_0�����H���źy�����sͶ���'L�-�[�
�����k��d����gKNy�I��#B��N��Ի$����g���6��R�>�-r���jښj3v��dƲrf���R��{'QP$IQ����J�'��e30�^W`tK@�y�F+Gj5�E;����-�7�)�^R��;�q��O����7M�[fD�[[7��<Ox��OTg�߻�lS���w#`�� 7Gh`0�~ ��T9R�h�%�eM��Q�uېe���EBuܹf̰���~����'ڪ�ô���v���2̻���� �+��U5�`�ڬAv~#���ʠ�SD̎/	Y�P�T�~R���jZd '�Ea�s�v�J���7�)�.^�=�5�H�n7&��+7)�D�e%�	m^	�9��
`-���5Ӂ~�N9�Jv�j��������I��)n$�R�����v��Uu�a�r�ә�?��\&6i|*�Z^�Y�ʍ<u*��������	�+L���H��c���t%�Ԓ��e�r�Z�O���2 ]Z�J�&	vL�<�I@��Tؕ�bg��܏݊���J�V�<j}&�\m���;
-*�sA��c=� �y�5lϱ����^0�ѕ.�O��H�{���3��3������b���˴(Je����qhC0s��:�<�[�p6�|�����\�ܻ�K2{�=������=���"
."�Ⱥ#I� �g��K�뼼3�h�*�?��N�aGḘ�2<m�:W�F6����4Ɵ�B㘻��3�i��Y�t3D�H_��J"Y��{@���
:Xf� pΟb�L������A�C�A�����7q ʜ���|�֠?��zUg�}�D2gs����z�G�T�k���eV�v[��y����4HW�gq�GD��sS�;X�ס�t�׽��ș��o��1�RC�C�i��_P����� NV�CȦ\�\q<��$��� ޵@oոr�Xٟ��+:���8)��T����;�5JƫO4��?{�9[�م93Aj��R�#��,�p>�rQ�rS%�Nf��_��i�*�5���