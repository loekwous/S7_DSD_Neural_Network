��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`wܷ(�D��Uݨ洅?�}R�$�� �ijI>R�B��e�h����``ǩ���1�C��1�%yA��H�ڜ�j�fKyUa��<
��N��8�Aª�wv �Z?$LC��a�ܰ.!1�z�r�0��l[�h��~+�7��˟.���H����~��U;�( �D!v�\�Nn��<�FŠ����aTA��P''q7�՗Ra���5������^2䣃��m�S~�-��\I�8�vx(���M�o�۟��9+t��[g@~���Q�WFJ?��j�Щfd$�;MP��Ҽ&�6)��*�}�������w�v�����#k�/��xj��I,r�	�z�@�����w��y��&���a_(�#�V�j��e��?%��$�hnk���-�/�=oZ�Q����Ei�26��}!�L�e-ۓ�,Y:��J�փ�Q��3��S����=N~@�:�6���WP�x��< �v|�TÇ9�$�H��H]K��(��N��^�����
(�|���k3]2�����Ѐ��ə�<�hc#ĩ:�2HG?�yb(_��c>a��7�(e��v�A�\�c���W��U�ta�[Y.��b# h<�{�MՉ��ʓ�c���?� rA�%8��|ܐEO������0�ڎ��a�Y/��]
��]��j#�J�ň���e�@䖂Zz$ �]�
R"������v&�w1��(Ňx*�ʈ�
7��X����#>�M�ӌ��ǳ��׊��&���:�a�Bɉz�vu���:"��P�p�t���[��z��ob1\�,nX�+��5��3~��=3���5��k�/�+�͏X2j�lq�;�ԁ�iX|&`�Ro��D����}?���մ���	�撫��h�AXܷ:����o�}�t�Hh�
O�#���~��طn�ع�&�oz�P�7���Ύҋ����S��_��@�f���j	�d��g�a��k7P��>��'N�m�%�P���9��k�0cc�7��a���rgpT�I�ΐ1���h>���y�����c��'�S�tO��,\�v^�}W����{8���v���Yp��ʛ�~W�f;9}9���pd	Z����{�Gf��/lb�3*���5^㶻<�P�9��'����Ѽ&�^�	��eO�v`f�ޮc�6/:̍���#Z��K�!�q|��]tx�D�cO
��G�f�l��-�	�:~m(Ɠi�p�+.��7`�.�A�I�d���8)�U���L� K�q��}����1
u"i�CVE|��I�&ƙo��P֏`M�.;��)����I���.P�5 O܇4H~1����4Z�5"3�U ~����a��+�me���u�9˨A)(������4�O�Q��|@n�"P�HW�`�[v�ب�����J�N?���&���å���m꣝)��H�G|���TVt�y��j��$��h���C���Ս���e �0��WZ(���N��j��e��Jc�|&	�f���k��I���JFL��o�Lx������d�s�����P���L���;�|����p��$���7��޶9�v�V,s����E�iw�<7G�d���+ҡ��=��f�˘p�aj�7���%�%5�?�r?2�L�$=�f�S	��_�ʊ���FIA	��'jÃ���K��q�߯�J�Y}�Zb81�RKra0N��!�����_g�"������e�'x���tq�_��E/AB.G�o��D����^ʢ�&g�mB�(7�p:U�ߛ[����	��:�[ʹz��Gvz��U��K!s:�8?ޖ���P��7��}�l��t�;�R#)��SȐ.��Q"�	:�T��~�n3�ݾ3�)��N@�1�ا5m�Ď�9$!���$s���@��(4�;�Vn���?�(?_4Ѯ(�2�:j��E��*�+�
���ziw:@b$����8��Sw�����&xySP�]��Jk�Y�)o�?*�?W�h�A����@�H��9d�uG�WD>S�_�WD�O���pC��\ �"�"�(~� V̸�hV�w��n�D��w�"��}���|�_�I����ڣF�͌0"۰�	������'T�`���t�\��kO/�
�^�'��Z�����W���bxh�+YQt#��b�1j?髩F�l!s�2����TH��ID��@�z�%��Z�h���qb�7����`��n� ��<D+�`C�+<�Ǭ:��:K�"�V�;_S�iB�p`�������֓�}�oNH����Is)�?�wF� ^$^��Y���	�%��Ñ`�������{&��<����� ��s�{��%��A'�k<_\(�ێ���n,��
�(׹Q�cȘ���e���S�Y��l���M�/U�B��=�Ӭ(��HQ����!Z�.��d��9²�!�t-@_�h�l�.U����n�C%<�B4�X%���"�q�xE���_�<=}�A�LA��F�<��X� �p��x�q��"��`�m��LI���h�{���>u]�'@��>���\��>�(�(��������cB��n�5��kq��m�i����m��u��
 ��>��Zh{'�L져�%��a��Yֆ�^�H���@�:�׭z�������Q��0r�xbC\.����r��� ��*���R��HN3C��F�u�}�_}� ��|C�BRm�ω��^G���C�_j���N�Z�c�^�!�0S����S��jzA�ɫσ��G���;[�^�f10q>QX�1͜c�4�s���=��|%�L���o��M;�=��
���Y%����ʸ���a���[T�<��C��?5lB�:�$+��㣆�La��a����>�
¶��%��Tus,͊��EHA�2��s˃N&1�kY��eK�þ=�{ՠpL����mU��ł��+r%K}����e	f	�j�7�u���g��ѹ[:�iN�~�/���7��'HHO�4=e:�ߴBw2��ϕ����qp��>��!P��$�:��٘����,C���t���R�O ,��{�j��TbeQ� �P�\t�u�h�'�tӏ��al\�j�����Z�@�Ɠ�v�����y��8SO���U':Y�1��^l�_)�r�ѷ�t;k��&`�$�{�GC��ɝ��c�K=IJtm��bx	yi��뎅�\���L"�t�j3�nIC�A��$�qyM,�|�E�B/������讶�Xߢ[¶�ʷa9���Qn2����2�2��Nuu�l�N>��37�W�㢋�;��8�ϘK��f<|��3z��OM̕w�����=A���/�(��P�I'ݾ�m�� '���&Cy^�+u�z�.Gn�ђ¤:�5���So�m����G���=��*.�B����sz��6��{����>k�����=`�6
�;o5gݶk	Y���P=�(���/!�"F�w�ޭ2x"�fUΖ}�<��=!]�_�wDB�d|���V	���kf��!�{v�ק�ƌ(���׽��w��\�(������Q{X��`O7 ��7�K�A���p���!���X�y�>�Q�{K�(l�1N?:+#����Ɍ�������1�r�%t�@P�Nn�� ~v�
�}��C��.Fe�}�b���0<�?�3�����Dy���I��a�ݼ�"��;!�c��i��ߢ)����$9{~L�m�|=V��$:�
����;�flv�U���"x�gٕ���8���3��7��^�%���-��d��5���X �.�O�%o:FB�����"#Ǔr�e%��e�N S�/.uc~��LMR\�O\
����E/�ۑ&�)	;N�<%��S�
�~ ��j���Ȥ��N$���OS�U�ŒN2�鱃̖Ń��,Y�v�����OiN��S�0�Ç�+~�}.rC�gS)��ÜD�Beu��x��X��i-�I� ��������#�Y@�%�ô����e�hws�fc�߈�k��Uv%�?��UGd�n���I:�?�@��@��>��-��W#��4�d���s6����"s��I�9�����q�2������YOۭ*��:>lai�:@pR��S�6��s�]H�� �be�h�i}ٟ�#�{s��%jX<����	T4r���KcΔ?�Nb�C���̿�dEۖ:�J�����a�AY�h�he.N��R`0Hs<��N�!�[�"s�/~W>���j�%HY��Z`7~���L�vx��x3�����VKY鳿JNJ��^n�°��(��G&��i�]<�~J�P���q\�(v�#����婭��N�6H�y��e��� �!�T�b3+U����1AD�s61jc?��^V@�2��{J�T���F��\,�ʲ.�����$v�4Ip5�u�lL� �1���]]_5{,��;0X��?��E��C���:���G����`�I�Qf>�D�7�.fm�d_Į�1̸�oX��}�Lq;������
Z�+y�uHw�\&{KT���y=�z!���&ן�C,��zY�	�%�:����s<p�k�&�i��&d��@4�·����&��sW�Aq�ĵ� ���l�G���X"�꤭`�����L ��!Q���ZZ�����е�&w�6]��:����@�_q�c��	��3�%�| ��?	W!&���(�%8Y7Qm�n��Z��I�Cq�U�1��1v4<܍6-N �;�3�>lPHղ/wh}�	镋��+%���s���
Swm����Ҽ��õ� �{ȭ�4��,|� jU��E,t�3T��e�CE����T< 2��1����C�/�����h��$�!�������t[w�C�I��'`�I����
^m�������j�ZBrI��x�4x�Yy���� �1���H��;��@w��ߟ�}��Q�lV�RJߖ3]������n�C_a��e�j8�v{���}�����{RK����r?ݼ���ƈ��:tB���'	��'f���RAp�%o-�b}v��)�����/��E���u�같E3TUs��q� �BS�������tA���L�p��G�n�G2���1]����� ���R��ژ��|쭊V<�<�����Z�H�͇�T�M�.�ݫ��4+��T�0�W���[\MBu�fd��^)�U)E�D c��7��b��&����:G?�@�w�����
�*��"�NU$�WSS�����H�2'XY�8(/��1z�����n�t�j��p��kږ-he�)+�$`��l��
4�V�a��SP����3�`3�JX?W��n��\�f�lRNz/^|#�iEiHLw:A��a�Lm5 k$f��WuuB����3�ֵ\����T!�B�H�Z������;���:thjPA�zY�.����|	uҌk�H�����fc]�:����B�.��挲Hi����S @$���J;��\��T���� ��{y�	��Ҝ)���F�a�,;r`�W���*+�o���L�!�ק��OQƶ���lg7��#��3�.�N��,Z�����*����tm��z/` Hѿ�Y�f�&;ɲ���Wq��{� �V�eG/�:8�X9I��W�B���*�3z.FKF�r̯.�L�cT����Bb����,Q.}��x��|���+
/:�u������"n:]S*�G�z����*���h� ,�XEEU�;��y6^�Av�6��E	:"<�J$�����z����g�H���xʅ��eog�IMU��h�o�hFl���$D��*�<�fżnL��y �9D�<t�?.�jet�C�GI�=��ht�������)��k��:]��Ĭ�I��"��)�W�N�蓂?\���X2Ȭp��   :s�� �Y�}d�`4��A�ʶ2�W"ZV�C����nM���l�A%���p_���a&�9���."ɻ��#��^I�&�B0����BEL�
2����Ʊ�$��x:�rOs��´h�Ͳϒ?(&+
�	� �t$��� ������n�Hy�u���W�1��4����}�5��%��2T��=���f��ݖ����<��� `3�*(���.#��h�	�x��֭���6���C2��m=�]��s�-�d�,���y=��� �^� ����#;�{�x��@�ly?������*0�C�Kza�p�B`1<��ϰ6-����*�	��7oo<.)8y83~������h�p�~�SjtG�6?ؽ)s���\�\��ן���	�����׶�I�i�U)f�����}2Vƛa��(���9^8�ׅ)v�k��p��&�C�6%}��L/5�w�+�Z#�J@Ӛ���!© ��i�8��eg�]>��������&�9�I3��@
ldI��|)�)w���k��"o�Ԟl���`�7{��-Ψ(��^�k��E�he����n�d�]�v��}r�8��^ @�W\�0
�19�0�!df�p@�"h2�����"_���#7�O�� ��q(<��C�5�OmR��=+7u�9J��Jx͡����5r�4� X%
`����0�w}��\ϴ�
45�!#�ug�r��\Q��=�z��-�y폡�٨B����P�RT�^^�1%X4Ɉ�x�� ��N�@C�IA���516��֔�PS��fM
�KEE�,�q�����wM^ ��[��A�u���k���:m��B��:Mk��:'d����m�pG̲��\�[>�����D?*m���޺��{�uW��ݧJv���o���bE���ݰc��$+�S篬-�M(�ʊ�f%.k��AG++�C�S��)�^�_���ިa��f�Z�>�����<;F�l��E��@�<��r:o��fg���7SY9I�qN��	�{��S��犂i�p�פ����=�Q$ &�W�S��p����,\��Y���"�������gхH�����]�PzT&Y��髄,ҘN��]R�ל�!�ReY����0eFm�D|�YA�Me%[W�QEg1Ka'A��|p+�X�W��e%�䐪$J�P��/��V4���6��r#��G�u�a7_I��23���),��{�FN	)���
�lAӁ�h����'Y%A+������!����~WƌDO,ʇ�^��ULHu��1^��R�⫉�R�G��JpҔĊ�V�؆�ϓw�" �L8����}fIт��9����'8��6��E�;߬� ���"��p�CX�Y��X7�5��(�=��	�/�q�/��'��E�e*_���A�O!���o�9j���WG��7M�w5W�CL���u�D{*W��ȤV02�]��4��^E��0��T��0-o�n՞!�w0dq�.���S�ܨ�ZA��b��#�t+�)�˭NU�U���C�@Z�T	j�YmY;>|�.�eAT	ac��r$�O ��+N#w��}[M�T�=�T�ż�Sڮ�w�H�;�On86�^���#�v����[���`N��Q���g���,hFyI�Mj��ˡ�3���.���t�rJ� ��|.���{6�h�I�g�`�a��`CPGzu�`s~��t9��B���V�K`����X����O���4�ʶ꺭�l�eߚG(YE�����Wm�Ͻ��Q��.�����)}��宬*6AgL8�J�{[�쾶zs��}o!]�Xt5��v�ZC�h[�D���R~@UZ[����bQÌ�x�|��G}��:��>-��V�}���`�A�WR������G3��g��ke0�,I�T����c��+${���4�j�ފ}X�C��z�Km�f���v��<�c3}�BEr�{~��Y�e��H	a��D*�����ftn�Y��9����:�B"�u:t�r� ��4�<�a�]�d#Cr��E�� �-�F���lT .�dR���]z:�u��u�#b����R���Uh�^u��89����u�m���'�콮��Z]Ho
�{p}�^�`��}5��
Y�� ����5��#5Ɨi@ӏYߞrj��9�)o|�ƾ��oei��Ԣ���B_۾�E��a��4'xX�VZ\��;����4���H7�G������K+sv��B�o��,8ȸ�;����${OD������`k�)&�8磺�/m���ܠ4�U@�ZR���ﴊf�L��,e��2�4\�G/S_���S���2��B5��*1�c� ]Vk�qkA���=/����֫�~_���}q�����K�u�M��N��j�ش�f����M+�]���mi�\���2fxSee�y!�=�F*��d��@��1��m����L7��?�(�LL1͘i'�з]?���uQ>ऍ�l�b�Z="5��"_�.y:"����2	j ��m`�;�|D9eռ8�\U[Z����+�}x-3�_�J�Qu�~���(��4:�������$���`\��J+V��ܠ3��R�5�Ffs �g��Y��X�BZ��$�?F��FI
UF%��PC7�m������F�/̰��X|�����8��ʞ�ŉ|���Η�xٿ�� ,�f��q1��*�e��v´)�y?�"���\VJ* �[);��׌%��g��;�BI[�wJJ�B�j��W)p������x�R��m~�V*������%�l�)�x(ߣއ���!�Y+H=N�j��ꩌD��^BQ�
yG���-A���N��� �=�J�1Y}�Ih�*�Pu��k����u�/fK�Ʒ��`O��iu���x�*H���]��9X]Z�Ѷ[,O{W&�Zr�Z�� �G�M�&F�pg���X��������&��X�az�D+� ��b�[I���d�r*IlF!��1 Pw��s|撛�;���Ψh,�)�R�ܞ�wdn\W�XἍA��j��3�N�i����m��!g�x�"�!�W(~���$�0�`4^
���k~�D�߉EN�^��,8̎m�]r���-�t@Gu�Q���2W�F���y���Z�LӾ�UA/e�� *3B,\��2a�Z��$�(s����W� �Φ1挰�/hAp���:ޥАu����t�f��+e �aX�q {��d�p#��?��ydu���+�SO��S��)��Q�Y�4�L��(/�	�h|b��g�c^�̝t�(����y���-�o�m+�_bir�H4�j� ��Sͺ�,���Ck�6�V������I��
�P�Ne?���U�z��K� ��8�1��#�\	*d������A�\^��w-��Y��*��օK ��ٞvށ(��B��]���,�s�p��B�Wk̆����p=G�t|��?�ٴ����ߥԎ���\���[@x���Xs���'՗2��ta�$eE�3ae1�J��`��9>�ډ�
�/���k㢐K3m�f��nH5n�SAO��m%�V���߇�N���4������%Kk۸����z��.�wx�RO���5�Jx
/��� m�<6��j-���&���I�߳�LK ��hV0���Z��a�l�D����;l[COe��hM��=k?�nn(��Qxy�(,���>6��o$���t���yp�;Fan���r�:�og�@� cɷn<y�˛��9@�����`m&O@�d�gDR��d�Q�p>#���]���Ǌ�2W�R�Ѭ���S���!�9�
���)�i��;ژ�ֽ��������8�ɴӊ�\�%��fd9H�}�������H���zTYD�6�_�(}l	/0;f���h1�7z|>��#3C~���n�~����	"����e�A�o`t��a� Ŕ��F6l�p93��>}�,C�#��s,��*_�s��E�<�WB��v�Ѹ��fG�s���Đ�,&<"9�1
\d�U�*B�kZݬA�3ǔ��&5��Z`qR�d���>6���楋�0pr�kή�R�(�p���^T-�zջ:���iH2������1q�A����
�cpb���ae)��)�Ib.�>��#���3'þ���C�U[ ��dTeE�	�V�4f,�I��R��ʴ�+�:�0+��j\V�i��I}���X����Ҙ	�s=z*��`��}�;�WK'h����G�(�-�BЀ�ymM]ܔ@�<�P��zKⵄbW�0B~5}l2��l��F)�y��LN��[���y&���cA�í��a��^ 0�[�'�9F�3�����9�Ǟ����p�O��6Q;���1�ia.]� �=�%��s(�R��ῤ�$��PPC�!�/��ź�p{�c��?N�L�1�Ǹ����-�[\���-sO_�"}�\�dލ�҅a��6��݀8$U���/�
�?��K��F2atI �h�]�TT;�1�R\���z�s�,j$��F���o?U�~����yuB����W9P��9�	r2��@��UZI�� ���7HJ�S��:s0u