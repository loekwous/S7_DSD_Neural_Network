��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�l�(���q�a��8`K�nz�w�V��� P�����"��l��p��2����}�iH��i�k��4'�����C�H-�%����c����ݮ�ƒ/L�o ��RD\���m#Ө���������tw��NA5b�7���ßS����2�+�X~듮K> �1p��M���%���|�8)�"���*q����E�x�-k��A��#����a 0�Ԗ~0Ghg�`,�i|v`����b���I���g �2|���KϦ�}U�+��t�qYBy"R�>D���tx܂�O3(�C�*U%f�[i��V�o���W�R�ѽ�	��Ǹ�L�8hG�]Ii��o�hk=t��zkC\V�P�0�{{M�^<	E�	��!G�I��E��/2T
�qd��HלgҚ������W�o/?Ґ���J|9�4��(:�zX	f���M_���j�)F���|�M+M+�D�j�eB=GF#�`FSF7�M��լ.|v��Ub��r[>?x��IOʕb�����5��X )�^k���q�����'̄�ThC|����Z�F)PjO�X�$4�G$sH~�u�c�p�������}y\V���Ծ!s�ċ��e7�p3)�c���H�V�,�+s����v��1$R�g���x��3	����tD���3E�[wI�P�t���5���#�8*`x�����=�m��e�)�B�gB�S\6��m��'<��#���bta2��[�9n gilZsk���8�S:SE��$P'j�������wM�X��]B�o[����j;^�&*�h��Hh��ł2=�#y����W�y�ʷ�Wd�7X�؋�KD�(gKJ�X�RS��{I��A�͏ЯoR���
�כa�p��G#nt{=���A	{b����m�p�^c=���Na�,�B��D��"��$��;���9y~4����nLܦT�G��'cُ6��8V�{������/3��x�۪���rZF�Fh?D��
U��!<K=.G4T��M��`Q��,�bYb�p�I'&��A�Ti��j~|$BR���&�Q�8~���EE �2Ym���kŔm�x�O�|`���(9 `��.��rD��UL[��ց����`�AK��o=���VL��{�F�"�&F�y�1u2*I��>�χ/�p��2��6F�O�B,aS���Z�����x�0��.(_2�#D�~/�Ђr����?�jڍ�;6	QK [5��=�˶w.)�Ȳ#�o�8���0����X+�C	�N��O�gHU���tA�2/��3w�
����	j@���~���B� � v�̻{�ʹA,��@��eȢ⌋�ߩa]ȾTy�� ����ܲ�@f:������J$������ aB�-��}>�����q<���)�b���^�i^�mN\�@���rz*�3��U��k쟽\c���� /ك�ޢ�0�2�~"j��sX6��p�=ߪCT	F���(���`���z�\A:�^���"H��U�ǘ�e��ٍk��L��>@rq�^���p�,=�tK�<��@_��>;���J�^�q>��2�XWj�A?A���z����d�X7rJ���_Q(��׋��/�Ty9��+�m>/���F�*�l�79Ѝ�T߹Pm��/��0��ަg)�m!w�D!����6�/�H��O�%gE{.�9�	��t�|�@�|]ޚ���dC%ڇMc,WB���Kiφ����83.<sm�ɀȑZ��e�q@0����ٮ-j��<������[���!��v�ae�x����aP��eo/���?��⾾)��;4���V�"s��E����4_������	Y�!`��e�,e� ��z��/�qR��?�v��>�jFU����M�3�wޯU)i��.��$O�Yq|�$\�4B9�1FF���%�5އ[�
5ؗW]�2ފ(��y]T)����z�Y��؍��IOUR�ת����"X�M�/v'E�4h����l&c�+�Й�����t]࿞zdk�ȑ��Ut���y?�N2�74�r�2VB���uږ�e���	��d�\y:KFW�fs�Oߢ]A�&������g:�3��p)mV�J���	4�����M�X?�P��pv6SŏA��4h���[I���bh�$���!tC)���Ml�E%�ɿ7�����J� ��`���븎^åM�?3U�?i�G��3 ���� D<�kvH�q�t�MO�6L�7+$�=p~洙�y��!)���|�y��1�ƚ���h�Z-��%�J����d�}�|�tu��P�c�os/���Bi�yA�.A�O�&�җRr�X��	^����7[	B��eRj�ͮ��G4w�cf@Y�>	�oM���Κs�I�}���ذ)E8;�����B� �0]��@c�}���<0ُ~��'^��Kh�����l��1��������-�:I��z5Xa����9 u-a0�0��u���I9�Kb0X`_q|��y�A��fO�����P2}ej�1O޾����&��O�3;\y.W�'(D�#�d\���7q	�Y5*�&omfcL�ńC���z�(� �ϒEQ��;�4x�����%)x�8��uk����7��kS��."|�4,Jy�V�܀Gv�D⁻�m�"�=�z×�!(��#�|���1 ��K{�b/U�Η���Hxg?0�/Zc�"}����3+�̩n��  �mv0��I�K�^��YWڣ幅<`�P
[�`J�nf�zo�l�����%���(naK� ������������(�I�}������|�A�'/l8L쟦� ц2��eRi�y�!�aH��]����1��P?�+�YM�k�:E��A:�W0����`i�?�ޝ�H�q�ͭ��+,_�d%�+�+���8��Qk��;<��Fn/os1�龎)#>��D��Kg
j���(�ߵ-�������5�-��x��[��F��ߔ?l�}�F�����_�R��K!����e�k�۶i�s�r�C�	H��Tբ)C�2�M��y磒�F��,��5Jm"=�������e.�^d�3%���ُS~Љ@�S��H�lԐ�d� ]3�I86g6��7n�J[�[���M�[|�d �z랰T��_��	�f?F�&7������þh���tۊ�{|��fDH����]Yy	�K:m����>|�2s�jLo�x���0�R��u(<��X-#�sM�"8�/hZ ��Ԁ����v������3ۄ���'����Od[�h��S�4t
s��be*��H�)�[RG��`��(Z^�t��U��(��#y�*r�����x��F����\_��Mdl�2d�܆����ɩ����N� ���D�=|�z��V��:i �e���]~$���d�㜷tccJZ�[]e��q9�������ĒZ��2O0��@G%8�g��!~�,�q�Jң�n��� }߲�������#\1d3t����?���b�-��h�%gܕT�Z�|�T�G�����R�WVc��%&o�����x���A���搨\s<�.o y\{��w~� �'�L.N`��Xl�R�p\²��0}��s���:�&������o\�����l��2Z� J\�߄E9�W�~G1�o[k֜�n蚶RO�4��׃�}D�xY��=�~J���&ld֫�ծY�9OѬ��"M�F�A �H%;C8��alcf�!�d�siq����}u��.ĳP��3b�A&��s��a���B��3�T�N�Ʈ(޼������1�����-���qg;���u��Mb��|C�9p�s���q�]�O�jK�mn��M��$�1�qf{�_Oȷz�֗��/v$���Z�6b7ĸ��Y0jpm��2�W�0�����&[�]�а0���)��^"]���W���׋�:Z�S;��9;���a֑��]����pq�	��O��f����&�i��Ҥ���S���$���ƒo8��RŸ��~k�tG߇��WÁ<Ld��G6�3�<���Ԝb��
�� �ӟY���_���Կ��⾊��C�OJ �Q^���=�U�䉥��b�-�C^n-!%&��Sw�-|���ˁ�I\�wX����I�ub~( �R���o����#�dy�`
RmY�1y��C�N�d>l�BG�|ɏ˖p�;u�f&���څ�1*9���TKڊ��>�9<�Mc�{�R_�Uyk;}�6���`�<Q�4�S�B|7
j̹�'�3*��ߚ�ċ6j��.�LԖG��lRps��d͗�a<��&q�O�\~��6���g�}ў�IQ��{a�N���i*�q7u��*��?ͬk(1A�Es���&؊p�HTK�V�e�l_�N(q�P�syz�%������l�gL�[[�=�(�������	���!F$�a��`{�t꿣Y|-z(�] �`X�%	"��j�����:�mٱ��yZ��^��_s�I�c��KQ-Hxqa3����j����VX��HaԀ�87l�?�4 ��&��I����vNg�����L	�e2��1�T����̶w���0�9�$ð���>P��uqx����Z�#�dG����� �UW%?q�$�܁oPϿ��%W�Y�*��ױ�r&��*�/��WU's�k�>���-��US��*X�`v$	M�`Y��9_(i�+{�~+�3p����I�8��	�@�U���B�-t&�g��*_Z(X���,h@�:;�$&����