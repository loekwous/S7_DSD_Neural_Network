��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`wHF�N�7�9�딩�iv�Q3��e>06����+�� ����Y+w�:���������hJ5[�\e,T,�'׋���0������<E�9��RA�0�Kn��wg,� �nC����>��f[�����]���0�I�X��!]�>����/�#��K�u�)9Ɉ�Ȧe�
��8��6%��*{�c�,n��� I�h�~�q���M��< #��Ǥ<},<bV���?MA<_~�%>G�#h��{(�~��à"L��2���ҙ�v:�6��H�M�a��|��TH���u��@�2���͖�ǵ���01"�0�Q7�6�b3���8���sߖ0@y����g���) �bjF��kd$U�d��m����^�Ob,��r�/��1��$v,ve���~od��&F�v<V�F��w�&��L��l�����<�7�3^�V1�K�a��!����[��U��I�`kɛ;��=�o���������@�����ss�M���Hc��^�����٣Y�0 ;�~\����
�����-��#��=ݗ����1y+���$e�CVva�E$7&�-��6�����$�
<�4Mj�)��f��"\�����x���{O+4p�e=>2�}�I�y���X�,�F��z7qQ_0)�b��������g�0�>�9�M5L-G�����ٓ+��l^�9�R(�4m3)'xu���Ǳ#�4��]�-�<�HI�6琗�Dd�ȑ6)ý�ę�fI�
�Hng�9u`x�3#*4n�8i�uC3�e��_�voW��R�K����צ.�g[���I�@�%$��)/̶'�&Gس�?f��+n����������#��7U^D�0�B�m��Q��*J�C8<׋;�B�����s�50ɹ��aCWO>̊�I�J����IM4Fq~�'��!�~�%b�G��.Sv�GH�9���.�!�#��q,�Ypܱ	�~H�����
�q�,=PT����Mp�r��۔%��x-V!p,"���Ǩm`m]��=2,N8�-�B�U�X�E?�O��8�����)u�x�u��ͼ�
vp1ߘ>����jHT��=g
�m�9��������-艙�l�k��i�� �h�������"~?Q)a�i�{���:���vK+�Ԙ�g�QN�-�<i�k��Gи��c`��El1���Nv�ez&���A����Y4C�N�^��<��=����R�٥Ul0̊�\Tk3���S�uߠ,.�O�,$�_��Ҩ8��vrYe��d
���1'�I5�=��6_��@k��~feϓy�HZ�V�(��9bt�_[�\#v������@q[�Pw*5^�ړ�=hpVd��ɧc�{�&۪p�Z�.Ê=�����L�8ɰ��ccܠL��b���|^���pP��^��
QȚ/ ���kp�!�ZKO*�ĉjİ��)�P>�ҖE��:�;�0~��F'ATlƬ[�]E�a�<���#�2�m�"K�x���F�6x�h<ʩ�J��9�>����O.�H/�s׌V�DI��O�~<���tM�㹊��KĘ�Fu:�>�?\�z�WYa�c�����Dcr���2��`\Νc��{�{�~P\v��!�[ 
�DL��u���fR ���U�qY��1�m|T�+��F�O)e�@�*;[��},�WUH�٥� #�	{ޙk]��>Ȋ^-@�y��G�^�@�4\ԐG����6��n�=|�����5�Ja�D���BX�i;?�Es Ք{�Q/��lb��߈O[��⤒����~O��X՜�i=E!�'S��Ǫа3�mc$Y86Pɉ-�n!E�$��Ϻ7�;�}|�#�����f�[tH�����r̫�h��(�~}��Y��{��*�bz�{�^[b��{����K��$#�UJD0����)4c�T�f%�m����:Sa��P%�^��B{Y|�BX�����j
���Ձj��j�Y�̪]�#��$~?@J�7]pMAm�nxm����B��O�RzbhD+�v�I���, �\"����dX�1=?Bg�f��ﻁ����W���)�,���"�؋>_n��D=M�F��Z#e�0l�yaC���O@�GmR��^aC�|i� �?#��>Nx}�h��kݿ�#�a�t��?�"jq���堯|X��DxgR9����m�/k��X�|[��2e���V�c�N$z��궄�so�C�� ,�B�
h3���=k:QX���ZxRz�!+O؎�F���d��ާ� �S�����߼�v�*�V����
���U���@�Ór��i`�������%�y�Zth���R�N3LrkS�9v h��+:�����F��̕Ġ�=�g���mBi��78W���7/�Jfz��ZZק�K�����dV&J�73��@6G%w�s�/�i�g���w��aBk/O��{����g����i���(�E ��/��/��X��_�X޲��h�v���2�ߖN$d�ν�0D�z��d'�c�
X�i��sw<�`�\sgX+�?����Q��}Ր�_������_���u�ɧ��8=�0���o����J{1n�Ӌ�M��n*�ğ��i���R�}���S�2��֚'��_[Z��e��������п	�7���
T��#LZ/yv
BNܞ�mhQ(�b� 򲳹�o����x�$p�d9) 
1|���5�0}2Y�R��o������(�Q7����=V=�4y=O�]tO���N�⠃��c�n�����	ЉY�-����K�ۀ�Y|��+n/3��H�i*R�Rx��Mѐm�H�dt4ʦ����:RT�'B����
��8Xت�>�8��7{���l�[�Q�A��ء�?4��mm�~�v��t���4�T{���"����#<W� �K1��7��K$�=��\&C�����"#��Z�X!���T��h��8=�t6a|u�����O�Yva�����.�8$Z��ël9��:+x�i޶/�)�Q�m�0Z����x5�H�szsQ͖zc���_�x�r���yܖ��CrFVR�{�kdI�g��U���Ca4V|�v�%�[v+Û�<[Z�ڰgk�pԐ F�`b�k!j%�/|׼S�9���l�q"�D潓��Ɨ��M��_,&lo�B��:���
a���3�Y���&��A���,p���f�\ ����1���q4�ac:��{�1>��\�p �*׀��)o��\��Xp�W�o�Љ�}��N�}D|q���A��Z�v`i\:�\����� @�QE��k;�̦c'$��	ߍ�!���&��+��䉃67�rUzJ���|=~'����^��c��D��2�/	H<w%�þa���򘙎׊qةt+8-Z%7�k%���)|�4&�?���z9����������`�p*٪��iޠ?x��(�� }欜(s��W�nQ|�Ь��zu~/��7�K��F�3�Ò�x�C�n��$$h��?���e�ۡ�`����s����#��G��^�	0]��Xn� �o��s���A�/������9�ӹ���b8��_w0
��O���i�m�WМ��1��T%��C鸴١Y��%}���$w$��I��w�l��K������^'�=�f��0z����44�҈��S�[ʆ�����*QCyť꣱��c׭�f�r������� �{�O�h��["����R��{�E0���*��O��"�_)T�����$9q\{�5��A���
��^)���ۡ�l=z�.;A|��x[<�p�z8�~�3$�Ά�E�[���ћA5¶Fp��S4��O�������a0��S����K�GZ�T_�ϛ�"ޛ��<��#��t+�*�XH���X:w�o�@�M�Nҹ�6xx��h�mm:f��E� ?(T4T���Y%��c�RRtdH�Wr�(�0�0<.V�&��1����{姆����W$AГ.�Bo�SQ!���N��=�"�FܤNN�I���o�b5�L�J��?��z�k��5����Rx���$Y;�PE���.�m<2I���e�\:��q�����BnV�!h�)y��'�B"`(Ȉ�O#s"�f_6FI�l8���nZu>����5~ج�Ѓ`�JI#��1�®D`�&�˅�K.�{��:�[��)�����e�����$�e�18o_d�����zÕXR�]vx�;,J�M�J���33ΎЍ�M{ '�Z9j��-���L�z����*]�x� ��]?P e�Fz/�7�?�	��l�����q������Yy|Ie_2���n��^S���o���`JQ׸~�������瘅�߅�$&��ò��AJ�/5�����; ��E�7X��D�6�pt(��%  ��}���
���^�]�,���Q��M�m��-'������!�e�����\N1�H��F���6#ә+�����b
_@n�k�$jR0��n��
�2��EZ0��`=�Z���>ӷ���w^����[�>c��k�����?��j�I���!\�!�G<C|Z"ժ��AB-������Zt6�V��"�}���9c�����l��4AA��}�P�8RK���0�B��*������#���O�d����s�wB���J�bb�#��{���bL{9��D�L�O����*\��
%xhi-	HNp
:�&�5��� o[=d@�\�؄�Q���6.OB�#��?Q�֧Է�s�
��gm�[{�ܮ��ǫ#pkƼN�1@������S�A.��j��Oxn��6����/Et�2��)E��=��X���*���;�x�����A�5HuQ�iU����3�!�)�A���â�1� ��v�*�^�X(�Q�RU���+�����t/(drYS�a.�=����])Ò��ᚅ�����5{V���ޯ#6�A�4��I���WX+���w�������M�H�|U�o����}�>s���Q�snB|�\�O7(a�,x;�z�	ef�m>�1}?,f�'v>�G��Qz/����0���PH��N�Cp�u�/�t�K ��J��a����w��z=p���֯C%����,^��'���Y�������y/ߌ�1;�n�6�
�s����v��D�������J��h��P,��d��9h����Q �&�.I�K�i&����A����^��h������b��N�V0
�`�n:#N��Tm
N �f��O� ��?n���)�$��åS�ocF=���ֆ�vt�ߞ~�1&������8���O^-]R����E���Ėó�G�!�<��S*���lig�"��):��黮�[U�	�[��0�����7G���1@K��
�N
��*&��tNd<r����P��@'q�pp[��ت2H�3��s`qMmzަ꠨^xo�m8��#��r^dVk�_Q���[��樯�i�Z{�G:'�ԪF48vi=�8�¸c�E6g���0��
p��2�\&�M�.A������@ܐ$��?&�8��˱�l\�>7�_m�M~jg\0�5��El����<��"��aI��6rq��\$x���"��1]��V|'��Q��1��P�ރ��w��9!_�{K��`��I5�#��ⱀ1�1у:J;���TA�h�m�ӌ��<t��J'\������9\�@�?����Y�ށ��8Ҧ��n�}mU��,,�A���f('i�HuK��y�0�p۶h�S�c�cJJ�6���!.'$��H�nzfmg M�N�;Q�����k ��`iO�����i�=�y�$��U�N!�>hH����;/?8(�ti���I�O�jQ�#{WG8hř�e�zH����/��&��ָ�P��6+�NT��˽���˥��R�5�Bqd/�+�����n�H1n������b��U#�n�g�",���o�蔢`�/Z�+.��ezrHt���
d�)�b��<�E��g�S �LJA�i�E�͆�=v}WƇ��ly�@)���4��m%L��o�I�<��M{B�
���NP	��PZ &b� ���؜�����<�~/@m�6�/<e�k�q�j�԰Ph)Y��y*�O�-O��T�8�ߕ��=�
�����C���t�E�/m{��7�
��W�"�$�?)fgqJG��O�y��r���������x()}'��}���h��!��V��8 �?i�j�0T�?1�?�c,�8�J�IR�)kG�Ou�0�O�m/�hN��u�r?�f���Wo�MH�-����[�}#�2�"a~���EB�%�x�����Ej�S�_s�b����}��V�Jg�3$ÀkaS��p�]�ȃ��\�K�i���bH�"�����8F��=����$8��H�a��1��.���
wcy�T�Mͥ)%~�_�':�^9w�� ��L�4�x'A��WV���!7����h�ܜ�iJO��@RC�
O&=U��)�	)SD���fnH�oe��7�w�J-B���hQ�"'�A�♩�Z�ru�ݾ��э�m��g�<�_�A�f=��>�QZ��(R���~�� ��������sĪ�
Q���g%�vU
K���E�#�ПF��F.������4ɒ�%m�O��k�x`a�,�����)S���ٽK+��UpX.Nc:�Ilq�?�F�2��9���}N�<6���/��gؓ2��XF:ǎ!���*�%~�R�b���@QnЫO���o�dD�O9��� ��Q�������c��|̕~Վ��x7d��x���ΒAlO�(�V��+݊�����,��֣/f�NJ;����=4�cv���܄Ϭ�A�%ؚ��*qʆ�٢Z�TQt��Kq`sJ\2)h����0D܆]���\b⊧�AK��	�3���Y�W�c!�m�|z�ӌ�6"Q�Zd�_r�n�{K����sw������	�c�4O�򙲖���(�h�2�GtspF1xI�\Y:���O����UO��UXI*�70�j�p�tN�1��S�S��x���;xB@��m�a,������{�Z�Df�[���� �r��H��'�Hv�M�rp�Uz<g�����OV���Ψ\��������Ϫ�+��p��0�����R�NA�ĜE�-���k҈�e�?����UF'�k�}\[��l��j��1y�Z��A������	֞�Y��ۼX�<&�Q��T�Ei�����.�5۝�RI��e9��u)W���4��ü�&=�.�ŘM�bшP֚u�5|/Ef�)/��`tt���r~h���Z����݈��= ���y���m.����_F�I��@alG��.<.���Z��z?�
�ݳSYf����(�=C*���.[q��JQ|�r�q���){ah;�Ԋ>�>I�k@ڽ�g�L���CF(a^��$��ոOio\8.wƝ��G�+�(��E��Rd�+Q��N`x@E�H����3��&��@��
��u9},ۿ��n~��b���u������z��+I9�[}���+���D�p�a_���LK���C�v������Z��>_p���� i_H���A{������ۇ�����!�4TWT6'rF���ĕr���/����G�q��B��S��Q�gj��t�������>W�y���ќf��"v�Y.�ld��4'�+������(�H��V�yb�A+]	��=�X�/*�񆪛-Ė��/.���A���Q�	�m���q���6�tNU�@� �m��a����������,��� Q);΍����)���ԝV�����31�L��#�u%`!�Q����e����P���SnGYO�UE
yyn����`��ڨ���YS��˕�q�j��]���ON���a
B�=XlA�s(LH�?ܿj�[��m�8.�?kz�G��X><�vv6.�踋�\���F]�X�����Z��:nR�(91g�0���/�"�G:��'H�#G�<(l�|6U6A��'цK�}��r�K����R�C���� ���0����2�X~Ǟ �������=JG���<���"m���}��a����%Chj��a�x=�а�q�R�1Y���ѓ03�m/7��q�駥g�O�ǭCD���S�<�>�2��y8�%q
�M��V��Ǚ�^��E�������PL��n5���qڐ�(u&cx��6޶���P����i`<��-�.@��
�e�s��PߛŁ��GP�. jH�9�t>��
�����H�_�����b�s�׶��W���=
 �}mW?ۍ�K5��p� ��.�K�w�Y��)�/�����pB��M-8���;���d��H�Ċ�ڗ�N9��5��No����H�'П��u�9!����o��5�z����!��kv6�e=)P5\�+Z�����?7�,P�7�֟Oz�˙� �F��YHN�!���r(k��ٓ����4�j�[赍(�LgcabD�"N|̭������s\�IC����u�=dMͳ��B߷A=��iP>9�!c�+�K�T�-R�z*v%*<=�%�Ǌ����t����87��,@h;&��Ӑ�zlV����,��
_P0�ɽ'�O�:cG�m��ط�T���?a��@�xq���l"��M�x�'��͔�<�{N#�lXi�����
��YA�w��7�-��K9Ah�
�$Ä�:��Jls��_�L*���]�P�)k�}�s�bߊ�[v�;F�p�x#<�Y�4M�� D�߄i<�W�\d3*�P���N©�Szn���lI&I `�-͝E����ڽG��+xA�*W�lD�)�}�I!/Q����Csũj0�x��T��J�G-F��I�"%����$?t�,A��;���.r�b�'��v�����q{М^����*d��Zy��6 RE��K���m��uذ>�v�2�tj����`}�5���B������n�s�L�r��͈�&FS�ȩ�ghҀ�ygsʁ)�F�иƱ��ZdT����2�������7d��in&�L�a������Tt�t��PI�g�?�۴^�<��ݐ�`FO>'����dSSt"�I!�3��)C28���873o�n��:O�=d&%�;��>���jl|����a����j�^+�5�ji�w4BC�_�T��G m�?��>W����%��-W.3�IϬ��VE����������wX��. H������;<�U��U�"�	��o�3��y?��c��<
|�d����W� ��o6Ov� g�]�� ,9WGY�f�T��+�ӟ��1��[;&�gm��K��ʂ��ǭ�]�o:��r逊����,�����3(l�Iq��֦k�zQ�|�λk9�E�6���Q��gF���S�������#�_��^ς�`���!v�.J��K4oL����A�܋�X��'�lu�2��B���lXo@b�"R[[#)0�m5���ho�P<�_���f��])��M׎!�5����%������`I���LÚ��zv��VFُ!�x��7�Œq6�[&S��+.�����c��8�	3��]�P*@@�,�S�x7_؃%_���+u��� �"�*�<���2��3��ܙ̝.�����g8�u-�bQ!-9 Q�\	Z�� cK�=�[��u)v�L8$��Z"���4f?3t����g�mz����X:od{]36����\oEH�jx8�%� -q��4�hM\YS��O��/���!�Ӧ�j3A�:𐱲�a5%�S�N1�`P�� GIat��o�p�-��a�ߝE�M;BQ3�;���M:F�p#?�6,1��Ф���`e�(r}w��/���&*:�H�����7���i�:ofp5�T�L�&N�Z2���? u!V�{8�z�$��os���Aʮ�����鵶p�U@��yǙ�����G:�k�ҍB��;�7��5��q)�6��
k4I�G�F�����z;j��[Ԫ��k� �,���dܾ���fGk��M��-x�UX~uIH�W�K���8e�l��ʈH����?b��k�ʫ���<קV���}ƂPM����s��.�S~�tva�=�wet���+q~Q���}�]�+܎��O�D̛�p�Tf���r���#K"��9QA���gZo|w�h�m���xzR�g^�ǁo,���z��V�:9���,�1�����R��I���<�;�����+<��4>�Jh>�9��L�:�7�1��ٕ��ؐt��m#Uhn$��C�)��m�4s�|���4]�7�h���ʿ����wI�T`@{����noa�!���҄�T�����!��F���l
8>V�Q��:� 4��A��V�/�Y�Bp\���t�`�Xv Q�-�g��ML�����6z�is�6��p ��*]�
vX���m����^�R"e��L�F��ì�JU*��K�3�&�6n�z�R��R�@l�4�}g7K���9@/:2��eu�Wq�S�;_�ttA�M��"��z��{�u�N����K��X���t��y/�L
){�.�bۑ��_I�t|�T%O"��V��i�q|�e�v@_z�7�¡�ڢ>M�|�̃$���yV|�	Γ��{>0k�̓Y|�j��;�_���h�%�-^2CҜ8������4?���Ɣx|���Y	��bC��i3*��2��5�m�ҟ���e��T�q�rnm&�3=E��.,�y��\Ә�"b�qX����D�|p��.�57G�27V+j5�Γ��z�r^(�n�9�}�jV]�2��|q�E��l�{�԰>>�϶W/�u�'s%���g��H.�YAɄ6�!�hr.b~�r��w��ڡw�o��.�*���A��h��������LK��U��S��i6>Z�E�T-���
����=���aխ:�p��WnѰQ�F����S�l3ؗWu�
#�o�����t���90��R�sg?�����v'�lJ�s:�Ob��agz���_��j�^����S�b�'�N6��3�*)�w!���5�,����6P��$˦�+aٴ����6�}[n�
J��5�Ы�u
9�;�ot<<�i���d'�J�S�E���hn���})+��*<��v�-��Gc��SV�[���l����_Z=jH���u6+He-w�߻�h�ۦb�%2T�I)�������[g>	�JBu�C�����k>�)��Ngn��: 
�h���H�<[��Fԉ�E{�YF7����A+�����x�:]��K�Γ��0������Ɔn*a%������ķ2a�2cj8D��\ӥ�����j���g��F�r��d�6v�__-�S��U �,��>�\�[
_�]ݝ>j����>��NŘ�}3v�6%�s-�w\a��*iSp���}o���f�;Y�Kj�W��5�y>�s�4m��U݌U�5�0��a��_�+WG�ҍ�<�b�N�З�'�Y�*�A8N����w���)(JO�w�fR����I��G�6��M�Ѱ�9J��)U�$�D��IT ҭ�F %�������F������ӭ�C��T�[�C�;~y��\��x,��}�.u�GF�t��/S��e���$ـ��7�/��>r\.u��xc��"դ�7-��I�x:i�j|�!�x����c�3ӹ�촬(�6F����>�\��Z�0����z���̼�r#��:�<ײ���|ǟJ�ll����þu�L���cd+��t�~��GXY�i4:�5�_�?֕T��:�5{�6t��+�k���BH&�Ų�ɕ�I�T-� yaf��ˡp ���o�tP\}�����c�
J�9^�g���|�2U�l�	d��g;�2G]�� �4�kjATMŤaVk,!�.��
r��8�����?�B�b.)�RKv'�Ȱ�!��^/]�l���|�[�X�EU��lcs�I�3�5I��g�
�����=@W��j�婿�����E�k�Q�3��v��8n�\�^�I����6n�����瓧�_�wt;:��z,M��~p
��R(�*��a�*�����/ż�����^���`O�K�`� \2%.�M��2�8A~k$����㰎��ѳ�5�e�y�X,Uc?Tz})�>��`6�!���:��Λ5�-�E����ݖe��B'Dr�����.�;�;��<yrևƽ�t��tG����:�Jķ�|�t���Y�:Ty߳��!�w�Xf�y{�ڄ\�M#nȑ����^��Ĵ�@b䑪w��w�AծP�x�������<��B�
�>�8�C�����L�H���q�ƀ�����H�;��j*�U���MR�[�tL�ibs�䂘�b��-Yrp��D���a�*D��B�I,��n/O ��DX����eOR�lvЉ����X{��-���q����fս�Kw�#5�܀�ۉ���M��9�5���!�Pٲ�L�9x�#�� �����Z+�"EPBސ��(���-C���J���}�@�O����č� ���8@���?�=�V�t�b&�~ES�N]���T��u<n�-ڃ��BC.��(��yf%q�3@�2S���]j˳}��H��w�Y�L��p��j�sŮ��Ѐړ3F?~���d�6e���se�<B�A��J�~��W��J���5'�REQ��C' ��2���rs�T0��m�"�쩃z��Ц��^+�7y��T�-�@~ℰ�t�*�(�G ÂU�@$�N���A��,��;���M���n�Dv�.��3�"M�h C��������	�A���s�D�򾜢�Ϳ6~[y%�ۖ�V�d��d���*�} ��	L�O��}h{D:ℨjI�}���g�q讕)���4�w;�����Ω4lwۮ�
&��ڨAJ[ȞT��-G6�+R�������=���ƒĂƿ�xp�����0�U�A��G7{X���w�Vn��H�E���0V�f���İ0�&���+V˦���m�����C�~~��6��l�7�6r������H�W�=��~��P���[���["�>��m_"�`����Տ�`��M�ء]���XCc��ݠ�ٖ����*�|�q���er�q��ڥC��w���Myt8>N�J��� iJzy���W��]��W�U�C���`��Ŋ�P�5U��a�5au��̀�I����,6�(O�W�Ex^-�c�o��?�ży���Lj��a/1��gD�^X���|�#���DX�-�;*�B�e��\�/���/v���Ùî�J��ߎ���¸"��f��S�F��}�<�n�S��37!F1w��yӸ�������'v�ܾ�U����So���U����06���{�U�]z�dc4=Ϲ+��8�3���v��ű/0���� ;�NQ<��6�&�n%� ��g9�=GHo\�\���F��+b�9ꨞ/��S4��*�-�%�j����#Ѻ���`�[n�I+f�/R.U0Z�����`�+п���6Tp�W�������ߜ棰�.<J�1斧r�ۦ)8�ľ�3
�&ػ.4��'|�Fh��]h��x0@FD�]�:�Q�����	p��/�U��GX��
�A|l��X�d�yMX
�~�_��PG���|Dv�(��`�6�Sϥ��N+Ğ�ѻ�����v~(�"r�ѧ� $��´�����[���x?SBk�."l �����i����`�q6%8ԃ����p�U.�g'��6s�)�dD���J�0YE!c��,�/��������u�
ϓ[��gF��RC�wr6�9# o��vK��ϝ�G5�㸘��t�'� n���ok*�L�zu�>���ï1�����}��F���P��>�����I$C�R~/muż�g�;�5�:H�MJ��1� �nY6�0o�њ�ӵ�װ$`�y� o>FD�ǿo��X��F�K��ݽ$��3�7e�W��]v%t����R����FLb�%L͑󿖹��i�r�#4�{�����OW^H�v��-Np7�6�3�!��ׇ�������;�b�5?�w��%g���Itk����V�ЖW���=ca-�[�	�SF���,� ��(��xn�R����eKh��8fU�-�X��H�Iy����;Ľ"�%��8M����i�6aT��ͭ0)�ӄ,�'%L�-��%�[��W��g��F�w�8��'��XDZ8�\�J0v��ZA�n�+��9��/6U�]�kT4r�J�+�	�`��R�׏?��I3��u��Rq�U�Sn�B��~����y2w��W]B ���E���c@N>75�g�iP|,V�Wl�����*��� Z��Z����#4S��Q@r�e�\���](���`�Q P7��%,G~��L�_�t�GGp�;M���!x����� j�o�|�t��V֙^�z)Ĥ����9ӊ��%����_M|�J�cy:2ݣ�h�z��[q�3�\8�ρ��u���,8���S�>�ţ5�m�uǛ���NQ��l��e3L�)������3�^s��Z���`Eݓx�{�\���1� z%}�iK%����e�d�6���B���w�ω��ɔ�-�9#Ţ���4�
P�kV�M\2�8�����3xB����̊�G
�V�L-�LI�ah��*����$qg!r��ѕ͏�@}u���"��I���_2���z��Q��M�U�ez���fk�j_��,�<�Þ���ګ�W.7>ꈆ7�ۆ�l-�����N1_�cK���O;�-���-��]�+��3(�eg��V��)�`�@�?	��抛���
�nC�(s��&>��}$��8�%Fޖ�j6T����߫�^3��C�.�ŧUq �"��ʣ��C�?kIw���|�8N<�V�%��7T,F,��yͬ�E>�`8��(lF:b$��=��w�V���8f�y���a/�C���r��H�/^�f�@�s��F̰ �I��n\_�������@�F��O��w��;M�IT+T��(c�{�s=��+u ��}ؒ�^m����'_�F���>�����Kњ�{N^�׭�����t��ܓ�}�P�P���JjZ�J���p�DU�1,���Wz�7�Ź��{����P��\8ܴ)���q�n9.��A�Ô߶��	sH���KY��ෘ|\��\R�7�U W��V�&rˁL:�N8�b�!��ʷ�ʳ[9n)�}ekMC����r���Q�!%9B*����`����׏QK�<ϳ�"��H��Ef�M���~Ucg&�&�r����$�~rp|�5�l��QYښ��<�dF0!4V�<ٿ�`�s��fN�"i
Ģ	_}���b�z�L�l���I[~~e	Zd��*)��xe������ud%4!O՞�e�F֒��t`��b��|)2�E�՗�O��c�:n,���(�5��\��X4�����OWh�u�N!�G�j������*��cD�G��uo[ ڃ�O܎L��<��p��+��$�A�Z��ᐣ�g�%�G]��W�'�D��k_K���#�W�<G�������{/�b����`���ޚ
���F���XR)HRdI������y��W�E(�R����o��c�T1b0b��b�kO��I��1����o�������֛L6��
}����>�r�w{��/����38ه�id�`�rx�w�L<B([�.��.S8&��~��Λ{��*)��"T�n�D�2��޾O�G��1�zh�� ���.�2��Ly2�� D��Ϥ��	 �5��e��ө:�fw��8�k�>=���7�+.v��؏gCW�����|��u�V�A'`WS}��5C!�l�����!����XX���fPer�x1���7D���sO��6TaO��p%�0�ϴÙ���:�Ŭ-m$�S���'�"O+��nҏ�D��z�\1`�v���bF~���u����P�?Ľ+�$�uwz���O���k��<�gl��:��oB`�!�m W��:�Z㶐�/{g@~��bt�� �g����;P;<s+~��$��?��J}]��k�PR!яj[0�1q�]�0�ӄf~$&�<�
B�i�������;mb<S��9��.�F���k���=&���Ӝ����'7;�&�ۻv,�ĝOڤ��;3���տ���_2T�K�,��4C'��.H/e�7�4G�"�\q��4x�Q-Ȗ-�X��1����E��J>��9�8�sT�d���fNn���,d�-p��a�v9+�`oqa�:v�X��֎N}�$G�7Q�|Ȋ,�L`rZg'x5��9��� ���]���K*��Ŕ$����jg=�"��f�;�����g_��gq��k`L9�a��=����H�Ag���P�y\e�ۗ�-�������6yJU|�/%� �D�Juf x�C�豔/B'��ʾ$����&(�Ko1�`��R2/�A�'�7Ka�_��n�۞�u�~8����܏|0��{��wUnF��P�s��b*�(��/�Ms��_��tJ��Yv;�N��ιE*��t�`�{��ՙU3+@/5	d}G��:.u��p+���`j����ejz��FN%�K
73)�u:7��k�h,����+c���?��Nx��-;Uh��>J�it�U�u*}���s�����'���7����a�o�Ok҉xd=+h�������\V�G� ��
�S�͑�{���$����g>l�@��]>�J0�Y���/6��0�
HO�_tPZ�,�YL����,�|:�Fǜ�P�j��pM���|v�*��G,6�³[|B���t٪����rH��;���~�;�9� �#��l��KL��J6���o*�]�����>	���ӫ.��v1��\�7��p��=��/�F��0ف�Z]tM�P?{�8�E=�Iٞ�����	gF�Վ�_�������c�W����OWz6�lw�f�,u6X�)�#E�����m�e��x"h���C�} �sԤ�
%���xF}s"qm逋��t�+2�h@�A���w\�J��JY�rfp�9�9�ٽ	��#�}%��4|ґo�!�b���TO2��9z�r	D���Wm�s75w����'�;v��]�/