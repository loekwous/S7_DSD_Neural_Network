��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w�6V�%{����"�`�-=@�o�� �ٗ1����E��).� �=�R.��o�Ӊ�/�~>�B�o�V�#v�qu�oB�{�w���J�W�.�1�np�ߍ?1�Z��V��aR�q�Y��a��;�Z�����G�uN���/O6�L�QF�\Q�����j�M�&�MA���E���	���ZfG��Q��iH	��p�li3�iL*�̫��ҙ4�X`>Q�9ߧ��r�"Tza086z1�b����+1~O�S���u>�:�"���
H�jY&ݱ�

k��r�c/�����:I�ئ62�j���!(]e⚴��ej��:פ:~&L���l�Fox�<bt�x�Μ�`l$l�A��8\�Ni�T���Ѩ��z�d�!�paEFN�`��H�}�9�+&e�=�F�>\5E,v�iɄ�}����c�P�Q�Hu|��U4[&���k�[�F5�C=d��Q]鸻oQ�>��9 ��ȃh��}c� �ю&R��P�p�f�A�[S@_ �T�8&[���I)c�Q7v@�8���ɥ�>����}�aH�o�k�A���3/�m.T�k5�c��;څ`�ʆ�PD�9Q��l�|�����)��js�o��BN����_z��q�MZ"ϗ���R��I:�L��77.�c=O_��@��H��Fo����U�����V�(���N�)��/���G�( 2$1|���\V�E,�N��l\���薌��F�Z^Ndm�ƋWs�'1�E��)�@��x����7�ql3�QUDt����|9���ϟ�U}����(u6�y�;5G����|?�K��������Bz����3��(�n��ν��<�r�q�Y��N�ƃDQ���"�w#r+f�Wn	��B, � 4��Pȟɘm����>d���n�x��o4�M��I�O���&W'�Je�kk�o�#�#���Cx�s�-�B_�k�1���DЧ����n��$����^��h��֍}ٍp��O��p�*_<�*��yݴg��h��Dl�*5�	N����ڭ�{'����|=�.&BC7���X�
xE�;<9{�'VN��>#%��֤+kv�c�W]�,/-���,��o�v���m�u��F��jrߩ^���
	+ۣ������b�m�I$�U��dX}h$"_)b2"��՚{x[G�����,P�O��/&�Q�j	�G-��A������c��oў .�-^�7䰯&�B#�^I��q��Rx}�#�I��h��x�Xؗ�~i��"�$�hcv�1M���!���ģ��	ED���m1��/�����ەu�� $��*�~Ǯ����k���bP
����۞�H�iq�<nI|K�d<0�X�-Ba��)�˝�ڶ5��H«R�F��u�^ŔEW$G�\��M�<�C-2k�qɘvPN����3/6 �`~��Z=��)+k�@1fX��}Tx�P�$G\�2�j<V$��P�=��࿗.�Pj�Jx����-c�(d�"��{#$�]���|�B��c1�7����D�9���IY��a��/����8h��9�-MN����K��72�ӊ���#s�k�k_�#���M0�Z��S���<�W��!�ͽ���B2��f�`Ip���? GM 4�ߟjYSq�{Kg��.��5�[Fc�����Ϫi ��%[��E}!�%?U���X?L��#њ�N�K>z��Iӱƿ���S�(���NS\���d3����ӈ1?���7D�ƽN�za���R��YQ|N��65]���z#{gD/6�,�Xt��9�o�?,6m�6j#C�Q4	y.?`o�`�Y���k�a��Z�rLх�H��Tv��6��j��b��K��c/��?�;�[���Y�0PI{�.�y<��}�W7���䙻<�5L�o�8�����+3�#X��<N%J�73Ҙ㋊pf�.�U~cbD�K�����2
�gIu؏�t�{{3=Cv�c'KݕÞD���k�0��n3�K�eNuf7��m����R��fYvS[�v���.�;L�$������5�vjzV�}�� �\끾h=��T ��F�ν�c	ջz�Ao��5�y�˜r!�<P�4ta?X2�Y�׉����2ɦ�/\���\��Q�*_N��7�rk���)���yÎD=Nd O�N�l�tW
�I�zW��	Uq�����V(�U:�q�j����Us�.�;>�����W{/AΕ,b,�P@�c�w?@F���" \bw���9|����g1�N"2q�Ǟ+���G�m8���ã�WwqFU�t43�2:ܯ��}���*�`�g�p_�n�Żw<=�wt���@�Z���|�7��9+��4g�o7���[K�J�7f��Ok�vc*�N�D��-�I�[o��_����M�L��h�
�*8���.�g�;��T�3�4[rO�Rm���������ti����.����?J&� �q��j.�C��a�h�f�u��N��8����)�����+��oT�O?Yo���G��^l�Gs�GwgQa�0<�y���Q�vq�9���P&]�Q4L�j���75z{���1i��Ĝ���g��{��ZB]_��$�	c�D��J��p9ᬫ�%���K�o�]I6��E�ދ�����
tKP�R�?ڞ�m�u�~3f��r�8>�уA����?r�{�]�`��j�0�XRw
Up�?�$��X��L�t�S�w������l$�/W�l��{��_�"�%�H��뙅�	��%���P�����C�5�+�"�����L����_/�IڣF��b��Yr���03�'2����a�p�$L�p�Ov!i��W���~=�#���"\[)*.Rda���Q�<�}m�L��8<��l�ץ��yiW��E}��[D�Ƣ�.|L	�M1������w��:l?f�@y�� ���1]>x�4�yE�|z��v�{������J��G���R֡�=��TBE�`����y�)S�l������B���R�'�����.-v���0!^��Q���������רj�4"���Ŀ�Y�����!�!�J3����o�J�iJ/	i+Wx�M�����D�ϣ��$�������u��9��f�IOi��`�)���-8���KR�0(l��ʅr�/�T��Pw:}��HQk���R�5Ct�Ev�u܂���g�
��B�@5%2
��[A���G�Z)���:�dD�B���< ����.�=�1�G��NU�,���w�T�mq����.p�e�O]�H�w"8�h���{����&Q�H�מ
۫������\�P�=<�U�	���ji1���MdV�Q�++��`��e5�Ga�B��i�B�.
ƪ�+ �ʈR���t���y���� ͣ��q��HF�?Y%�F��,N��b�UK��z���[!YӢ���l~�I�j�l��mJҕ�a*6�u%���^�+[L["s�0��f��t7�SP�����Z�� ���Ϲ���C��5���ķ��<�8|�xq�4\Z~گ�;��R���w-³��1�c��_�Y_��k��qy������p ��Ձ⦄��|Y�}������$�oi��[\�MH���{��#
�����w� �?;l�-�*���=���mE�n�J�E�0�o&�gS
w��yRѸP�w���vsFWP3�&�������mQ �����	��*�����{@�H��+R5aX�����Qy����"�a�~�ɑ�LH����e�k��i�C ���6۲���&�T��_����v������\�,���0#4n��[��`�^��/�UܗQ	���g���h��љ�����:BQ�=��Ss棉���=�ko��|J��#���Wg�H���~}:��YF�oIK�j\�D�.C����.y �!ȶ�v�v}��40��?�-�!(f�-�����/�����m#X<�<�`l����)z>���cׇ��I{%���"����c����:�@�Y<�v_Ѫ�6������,eա��Ծ��`������"Ҩ� m6:%6B�ml� t�ɭ�nD�5�N�u+���^a�t���-	6yO��܃ �-=b��p��昿 �p&���p�,�-~S�7;H ��guC���E+ YGO!Q�p�+�� ���AeS��)���X�˙�AU����T�V��,�<Vn�/W���^���KN���s�0����0�ڹ�_�-�x$�y1�ǘ�_���'#��<���zu�.���J��V��̑{�ȠVE�ix�ڐ`-9 �T�����b���
;�,.�՟	s�6�t�f� Q2$]��[�ӹ�>ʮ�-��E�p�O)��q�6֚�3gx��ۥ0��ٛ��g M�.P��5�
�E�L�)���P�گ�#�_q��*J�%~0I�u�$��w����]��Kyf:/M}R�����&ƱT���>QѪڎ�����|�$�
��(���Ҕ����tI�?ń�ڣK4t��K�BU�<��)i�,���M�a��H@� �J5 ��ǥ�w@#cA����瞦�!{�R`��@�m~~�v;}��o0��l7=�%,��t�(��rK����߶4�S��:h5��+�����Xԏ�mR;b�qpS����[پqpv�;?`�pF���x�qY�����M�Fw{���
������{�c�9Gȼ�W+,<�O@��r�6d��9TCj��TX!�Ԫ�=l�Yx�Lf'�� N%*F�>+�`�� ��_0YcF�3ދ����˞���֕�1/n�9�:���y��/O�Dz��6�y����(� d�5yv�
r]awH��:���~�ZN�A"�3����2���4���Y��N�Q�/W�k;8Lk��.�ұ�.#}�y��TУ��.3;��E�Q� ۈ߀���V,���}>�t�[��R�Y�n��I���L.�w�u�5fBP���ER8-N�R@�#�V >�ᐬ�������X�_�'j�c�;�n�0E�3��'M`�!ҙX=ڔ�,lO�.�a���t�aa����y@�帓�!�����hKB0]���wv�Ϣ$'E˜����i�w�T�ׂ~L<������D������S����G�܆���9����@�7üfD�� � bݘ҆��|�V�%��s	�K-S��s���7h��R��'縊}��IF@L�@�Z"@���t�&�������C��oB�E�v?��S�rN0��:|U峟��sN���y�Lxx\��%��2��v����UDΧ��U8]d�O�� >�R�X*[
�#�-;x,y�k$�����Z�C�/a�:S�x��TCոp&�Ac��� *����И�~�J_l���$�K�D@\�#s?��Vו�g�n��?o��^ls�,O�I�Y�Q(�>�E�K/#��rQ��
��v��j�P�GN�t�i�J,H'��)r��� ���[�4\��D5��שZ�wY~�aJ�9P'}��a���n!�d��C*�y�#�AZS��	WS��*I,�V�ٟ~`��Cj�H���덅�=���d�͑�b���±;+mL@c�Ox2�>�"��(thz�f#���Q�u.����p`�q�M�u_$���g诺͸�V�͟�/wh�频��i���e��;?��1\�^�����A����5(����a�_�y�(Ŗ�DxG�|B������<����)����aFɦ	����|�������4�RKn�M=���^��$�%<Cט]�q���=W����q�tg��)��VL�c��,�|��2�w���b�R�#rP���FpM`.R�'��c*g�F@p��G�+�[t�%��d:�8�a$4gZ2A��3*�v9���}R�'����3��ث��^{w�s�R
�&���u�J4!dJ��;;KW\E��j�N�з�/��}T@�����J�U� ?9��G�,��㍔�/����9� ^+�E�Y�oi�E��aι<;別D.�'�U0���=���N�T-�	����*Dycl���ʤo5�ۯ`��������U�crO��+*Bix�a+���_ ��rGx�>Ae]�����,�7È,��$+B�j}"��ri6����y��7��F�z:A��c������ �2�D߱J��'��]��Vm
:-l�o�]�,��}����@9[j�фO�N�2_;v���t?lQ�M���x����~�K������I������/d�]VL�b!�!]�S���7��"˧�qV��ZN���
��F�d�34k��$=�]�bjhHdݪ���3_B�m��n��ܩ�P��SM�J�9	X0f;#�"�&'��p��X����:U5?a����/y���C`6�������\`�,)VwiM�jo����i�f&:�z�?2l�f�7F��Y����
]O�?�Li�q�rv��S����
v��o�
6I�qH�5�n�鯦vd�>u��2x�"���f�Q��炯���u���#Ɠ��Ƈ_��G�7������]#k�X��9�<������ų�[Q'�dV, �o[�.q��?P�c��"��z^����t:>K���ιܬ�uD�VF��B�+a���Sb�=ј�3������I�uq��]	��O�Q���p �v>��塶�d�mZ�0t����8q&��ӑ�-�7H���g1����\�r/��Ҳ^���q���v��.���k(2��p+���AKq��|�6n\�zQv�3!�ќ��IːS��߹Є���b��Q�|�4>\��-��Pr��V%H�o���φ;�q��D� ���w���9C����{M_��[(���؆�sB<�L�^��:��!�`�.�.(��m<���K�@N����e���ߔ%�OcU�ʘФsO!B+���Q2˻�z9��O����a�f�y-��O����c�����ӿ�#������d�~����q<GvKB|��-(�6,�z�3�e�Ē���p|���eoW9B�x�����(����X���9m��瀈kn�:J�����⭽s��䟇��;���\�r�m�_	K?ރ��)�"��o��F��[~m��H��=��L�r v� d=$�?���n�w���f���d�f{�dT�Lq�DP�hJ]!�1&H�_�GyU�,���W#���^<ي�ͺt�K�H$�L�@JT\?�b��o)ݳ+��v�?�\v$�	i]$��6��A�����1�$��v��f�jU6��=�]>�5���d����V�2�?�`Ҁ %���4KA���F�J�:otE�9�À�M�tU5��<�O|��3N{ۚ��w����^��fv`w�`:`�m3��	}��i���F�"�Z./A�q&�d#<3_mˈ�!����]a����Ӻ*��S5�(x]Dʛ��2�=��{������PiӗS�dXcN�)�Q�������孃<�;R^��B���G��gO/s��G��Og|	^���|G,�`�m�>��ܻ���!i+�U�&bH�< �b�Џ�$�G��-��|g�uЊ�i�D��<�����U�;�/AV׳\�Ւ}7+���81`&��߻*�5�g�):)��Xw�N��B&o-ڝ�$h�a��] �ړ+c�6Â]`2��e�IM��5-�������W���I����%�����{������vOi�)܉wUm��M!�'�,���I��8obx���10u�KM�7���Hۃx���� �= T
m� A<�0I"��8�O�1���MCz֘R.۴������΀OXPt�a��gL��Bs��[�&TR֨��C�[�n*�ݣa�+�d��Oin��]�fw���7��NЁ!�|(��������K_l�|a�kh�<�-X2�:G�OTl*eC��5���]��4!ʫq�_㬒���.��<���7v_,9��}�T�O6��RF�����S��z̑'S�p��F��ru�Ȯ}�*]ۘr��	ؖ��G�?�By�Xm�H�����t%v�{����yew��q�?9��2Ʃ���/ĪG�/�E[�c��<�L(��)���>���L�d��>���ż.��وum�>l���.`ᄑC�	q��A_����|i���6�Ou�����=+t뀒�8�Ͼ�YS���oL%b}N�� �l�M�x������*%t�*Ns��4�xnr����r��Q��T�Y�Wv�Z�����
�C��wf9�����%���t���jg9FZO)!f��PYu��7ۏi����r:��1!38rG��*�p��߭ ����a��������~���%S��� S.�jʅ�$�5R��`D�@D�,���w���j�̊�����(�V`;��'�3�9M)Z� ;�#��~�����t��r�Э8�ׯ�y�W<�E\Ѿ���r8׾���Q5���^~O���z�}���Hf���d���l�8��U������8%c�K�x�$�G��k��!ӭ.�C�8�bd�# ��a��u���C��X� �7����'#�*�!��0	#��7VZ@݂�Vp�b���as���j�OC���{ʴɥ�#�I� ����� p�m�0S�<f�y7�g-�pm1�gh&}�-�8�΅��>Gf���f���r�-s�'`%#��*'U��.3�ZLί�ci ��I#��Q��L���#�[M�F�_�=�0��t5}r4���UM�l����#�ԇ��N�N{_v�C$�$�C~�-��!�[�~$��/��� �WL���$��׊�t�c�n�3;�R>���w*Vs������r8)0٧�surB8J�C*�3+EZ�x������8�\�8y�����z�6J<�4T�ŗ���,kU�J
���Dx��eu�:��y`Z�����\�ݖ�'v��?p�X�Y��%F��Q�2/l��6��3����瘨0�nߵ"��J��go�����Q�����Õ�9�Q��tĺK�W��g��#:)�V$��RW���<V�F�,����Ytmk�Ҕ�|�^E� ��[������eZ/����1p���V���%2���7�O��e٠0�9i��+)��I<͟����G6j\��fr������������
���B�%��M���'y%)������-=��P�M�#�~X��j�lI�[&`�A���uh���}Ұ��T����G��*�n'��$;�뙄S@@�g���L��*�vZ���5���ئsF�,f������Q02V����ᘞF�@7�
T��ݶ��C��
L&��/�RK
迅<�aX7%��}�G,[�#�7������O��r��� ��}�������p��c�i�_��
��D���-��7�X�{���=�DR�W�<!�m1MG����61]W-�e
8o<�o���Id��W��x{9h������^�"����ļ�k7f�1P�<4'�>���r-��-=�V"��(��b�d^�D��!�ʟ�<��a��9�O@�q{��R		��%�K��?so��:�D��x�J�t�L�QeA���r�N�����d7R��y5�0C�K�w變�*{���^#�9�*Hh�N7��<�������&<�2�v}��v�f!��7a��A>î�G������5_Ƽ������\���1P'�,�_���za���k��u����i]#'������Ď@����e�z��F��}�nY�z4T�Se�rL��s�����"l�$��Mk���-\�1� H�%C�!�����t������%{c���|}��Ko�s�O�vʷ�gx��R��_:�?�����.�C@�^�LT� c�|��0V�α�Nw��\	�_���s�E�������co��v��,��d���1&�rE=��r�b���l��[v����������5O��n+,�%h0�/6�k� Zo��@cE�a_�ےL>e����0+�c-@��+���<ήJT7,R�,[b!Q�9w����Y�
�WV�/�t���͵L��IU���ȃw�pX�)��\��@�]bBV�d/h:8%������_�%TL��X�47x֏d̍Xw���l�]�|^n�`���Q?ɓ����[�(�I������aJ�Ǭ�eK���e����ڰ|�P���f+J86j&
����+O �R0�{�T���~*����h����y�8�.�Wt.v�U^E��1-N� Q	�t"Z{��xK���g��>J�.��X#a���^�6a���C��$�F+�ĝ`#�{�x����+D팋��&@��
c�������
نK vV���(%���X�Kb�7>JV�$�����ӳ}ؾ�;a��t�6-�;G�?�,�%f��<T%��+S@�1��.+�ڔYdiYgP��F�j.�i���\�a�r,�m�-�Z���y�d�����7�J�>�C�Z���GC�yz���>�/,�h��V����2���Mg��^�<���yuB�cJ@����D���c8�ў��/�G��E�W���t6l�Hk:�p>~���A,�9�?��M8��uP������餉N_$+6*��=��X:��&u^��{���nR?�}�I~��u�@[Ϸ��jXja��h)��T���,��&��N�v���K�g}S���ɵ�'4M�ܪ��B�#�]��R;�@m(E��{ԕG���n�)zNiI��sX$����)�"����?��'��b4_�t4o�7ɏ���7CAa�J�=S��#B�Bձ��Қ��_ƣc�KWZ�ꖱ��=��Z�\M[M���k��Zѯ3=47^��^�o�a
���Q����.��Y
*.����ԛ� ���=#땢��:*q*�>ԟm�iƴ(�PCQ�+��j��%nނ���j	(+,��������=��f�!!�~���0�ӥd2���E��kԷ��o8!��.�q�[}s�3��fd��{K�c�]7Ά�~-X�lWF�'�K&��]&�}y��Gt��Y o@��E3h9�Zc�F���������,��^���a��d��y5�M�	ξ��rv.�s��ʾ�\��k�p���2H�
��:�M3TՂy��`���9����l�Oe���M�Kޮ�g,o��ؙ���8�m�ՇJZ"'��A� �ib�_]<C��/�~X���H�����?XՔ�bM�dd��t}�1�vs�Z�y���>��Ep&Ԡ���ݝ����_�鑷f��r{s��C���̰Q�	iϰ�8Q�
�Rxx�]���,�Y¢Bk�����
P*��8� ���Lm.���e���`����]�"�.uU����\<�˥���x�{8����b�O����Xv���N��KW�~J�ͳl�����~}RB��+M|��5d�۽>	0�Ak�F8��A~���+Һ�Z0��q�r���x�W+,�ͻ�
~V�ݪ<�	,''��;�vS�P��`�����o�&��R����X�����y�,�X�v���^����m�4�藳�̫fj]�@��T"�w�	���6���4Va�������Ũ���H�8��')�X��?C�����r�<T ��$��0,�yW�193�K�FB?zNWP�ܱf�F��0�0=Cp?>�H�gUW�t#}L�B/��nS���p�8o�L��S4�-(﹬�l�f7��*S�QT�� �u��\��PW�٣�[_]s�:��.���oʏ�ir�,��6?:�KN����I�-�7�c���@q�����9�J���	i�A�;ĭK��:FU*�>�N �(%9�Z �j�����C��֭t$1#��m�ؿ�Z.죁��`��q�8o��?}�/{������g�)�f�/�Z#�hZ:;��;o�v��9,�I��?w^$���N�W�7�Kؖ@�i)�k<��9�n���rKkt�x��bۏK,Dj�H���y@&����%a ށ��_�!ܖ�F���d� �&V���n	�� tM��$��>A���8ǐ-~�Ut���UͼX��4v�aa�\]��!�( ����B&d�%��I:���u!�����_���i|��t0��e��}�������������.�$��JI���gdj1����r#)��L���1|�����k<�����͉ޘ��a�ZL'��qӴfQ��]J�����_T�T�[�Y!��!���KN`�K60��R����GT#brL����6jXOJ�n"3w��x�E2�Ֆ�?��h��%o�V�aZ��z��|�͖�qPAgWp"�,Xđ������`z��5�#�_�W����IU��(/��m�I��4FՀA�p��,��2gp�ꨩᑆo ���ђ���?�oಽ7AlN,��WI�[Q�0����d#�?ǲ�-��hI�D֠�f���r�l&�U�,鿠[�\����Ug{q��H�
Z#�eJ~�U��I���C���1���	�86?�<6.��D��f\!l��UG�?:Og�i�: ���<A�j�[ZP7s�I1�޲C�}�V�q���ȟD�a�o
�˰��pQ�'�8�q�@p�v�l�[8Y��]Q���v'N��`Z���?��X�)(6��
��(^0Ba�0�5$�^�;)&�1� ����#5�{R�x�����2��M�;��tw���e�a�pvQl̟�#K�����Dy5�%�J�` "�2sʓ�{�L�G{eb�2o���Q^'4��b�"�)d��!�N�j�hI��Tw]��p�(�[�Ù݆Eψ���O��%�jRTt��E�Z����t� Q@<`J	=�o}[�G+-�l���y���]G6; �4�Z�{��t��Sg[#u���iԳX�]�����j�1f�1����O���Zx[N��w��RpA-ay}��@mu�>��T�1�^��}J-���$�J���x$l���Ǜ������ә�Lp"�`{}��D�%�ҭ��0�Qv�!S�k��v^1���X��0aM�#?�q�
�!��^!��d��8��cI�mJ�O0�1�06G�����x^4ie���k[����n��Wr��Pjo!Λ�$D��b�ȣ��k��yS9�O ͏*�E�'����$԰�&��:~6V��?��0#��_ �6���ZLO���0D)�z�r3�����ߍ�N�������p�P�2n2*�6'�<aE����G'!ۦ����5_3����/�2>NkN������d*�T�����	m��Y��z�zj�aaQ~�ˆ�P aV�U�V4r��u���!�u�["{z�y�L_\(?�3��颪p�� �h���� ѵ��$������ %_(@�~D@bD�Il�&Zu��~Z��̏���������ӵ�wd�f.H����V�޽����;�N��4��n.f����q��u8�P�Fd$ڴ�r���]K���jHV�a���n����ⷀ�d,��G���Q4�~x~��V�֎A)y%���Q�~�����]rIjֽ�i5���d?;��T�*iH��'�k��GxeF�8_"�+d⚉J�����:]�s�Ek�u�}��!�9`)FV������Q�KXu�D_9�r۫��c��Fһy�������찑t�`�������27�BTRgO�N ��d��.�G3��.����4S�,���.r	4":8��"w��ᧃV�7�7x��r��0A �w�u 3��]�e`W�/n;o���y��S6����b�m�����3�K?��w�B�b�ޱq6�楙�\��r|}�����<n?��wQ'�4�e�kن���E�Xh��-Uf��r�Gd�_ufU��������N�	��8ϖO�R�x���O�`K�]�3$�C\��
��S<��'�O�[XK�b^�߂ycT�vŗ�\WN6��4W{�B�AfEþ7d���'���3f'[��Q[����&���1��/����-�I֊�)Iv����o��z
�D}~c�LW�4~�y�I�8uՍ��1���}7�3�EI)t
�̟�˃��jVZ�y�C�n2��5�Q�wߤ���4���#�~��L�y� �r<ő{Z�Lś��0@���Be0U3kΊ��ޥ��'`��Ռ��sq�����+x/w�L�,zKm+�"|�\�wo�V��R/�_�j�q;�T�!�t`X�4��H�@��f���y0o/�D!TwȆF�I��>�%N8����g����$�,�\D�7�]���yA�A���8��M�VB"�)��x�r2W�zb����g��[Ӄ1ˮ��s�M`�&��u`&YK?�1�F*u��]���HY� al��<��]7+�~(#x�?'R[7Y��=�_XjW2��>r�eeT�(����fE5=Ɗ��/h{DK�D[2XG�Α�H	��T��϶���hkLY�6���"uݻS$(�\*[�DJd��`[���G�K8�����8��w狵��5����0"O1Unt:C�ښ<s�HۧSO�ݔ,�Cӣ�f�����"��7��Ob��C�����ŊQA�d�PXF����K�]B���l."�w��AgO�멧�����n��*��Βb*u�g��s������Z�"q�Ȉ3�QN;����Ӕ�֛L�)��b-��>�X_!����'vz�6�Y|!��.���s��������2O��E�k���Տ+����cXL�
��.�ťX��`�1�j�)����^���~SVh�����S�4k�����`o��$t�������W��f]�g�²�G�c��������z��N�N���X2��6vuPD��r׬ �3���&?>�)����`G��@o�Ld��T����T���~�W�5���[������J��x�]�Nk�ci]�dK�Y��c��x�SOٍ9��h �F�
fL�X1�-�8��� Y������=c>d���i7�r��a�L����c�g�w*��[>µ��:�]T�gL�6�B��O��~dYբJ$���G�@��'㍇��{�_K�{�9w��j�3T���s@z�w^X''�<�7J��"��}W0��ۈ���(|ʓ�O�P��M���>45N©�Zr!�0��;�&�S�=v(��9u��ν�{�&B��Rw����,��ڟ�
M����p?yF܏���
��[�e�.ܥ�ul��q=l�s�l�n&�ي&�H����� ���bي�c�X�7��C.(����[��b�kŤ/�������)����̘�S0����Ab�-Rf�_������~,o����"YAUSژ`2ȫ������rQ�0�z˟S|�r'&5�x5�K�o@��"��5�����}�����S�U1z�J�叶%9.*�����|�����?d�8�aR`�m��.�!�'��"�d�Z?�f�M���ߟh|������2�O�>�5�ȝ��@ǯÐQ��\Ô��|! �!X���*5Q�&mh���K�aH����;���� ���vS1�j0�]�B�[�C����_��{gE[D�5��%��m�i�I�JL���J�`9��t�]H�U�l��w��
��������=����_�W�D�O����(�??K�'|*�@�?=+�3,��d���L�h��ݐi��t����ܼ�B�+�#~�
�?z?Xֺ��$�>�}:�f�׋L��!>1��s�C��3�j�,y�P��z��|"�3�z� #�l�o�/���:���^|t��-NA��[�C����@j"�Ou6ᖋ^ K,�7�d���n�ŐN�T��A7�Kv��4D�n����"1���[7���үě9�����(�h鷌�4Y#4�$���d{��z^L���)���6u���li�¨����E�6j��m�v�c9���������Af������C�fκ��ԛE�����n��[�i�n��Z{rq�6�G �)�U<��M�_wFe�.,�9sj�;E�1�`5FR�<g4�u9W>�Q���dlc8�N�:��2�?�\K~���R����4M�&t�݊��A1 ^U�^��ų;c���ʹtz`]������ĸ��?5�I`jI!�vQ��.qQ�97�Po���T���T����g�9>E�\�p�dWB�Y���Ɵ;�j,1���VK�u]����2�>��.x�0pw��i�|��k�M
���
��7�[W����PK�Ͳ���7n�f=*��W�p-�U�L���)!�kGö��Q!J���i%ޖ�P��Ԭ$�&*��b�X��'��X�k���/����W����~4�b��^��m{jL�����ט ;�RH��k�y��R2���6&u�\ ΁�"����TE(h�*�-8�"�ص���Cigء���5��]�_/簈��qz��pnKUW�4DQT�S%mh`�>��t�v3�f���,����	􊞇�s� oe�p�-Gi��0p�Tn�X T&���dY� ���3A�RC�Ʀw�u:!a�����=���^nHV��y�����ի(pɶ�����o��k�ߟ�c���7�����ǽpc�R�cM��%��:�hƔ6���ˏ[�\�LB�F-�ĝ�0臟@�H��	�J2��8���b?�&�R���[�;t�9 ��aCY�4��$s3	�}/�� U���7J�B����)��B�߷QÛz�RQD7#�?�΅t��:Kd��3�V��	&�<-�1P�:c��Lʭw�ͅ��d��_Hw���(��x�2r�o��7׹��ԃ��!�b��F��ڏ��x1��h����I<���bh{v��[%����%@^N�D�=�N�컎��2�35.�t��x�~����h�HGJ�s��qU_E�<Z[��� �I(�X���w@�p���h���gp��A/����L��K��|��7�	�x7c��*�$���4��:�U�hyG,������A�a��w
���"�*v����H��P����+�`��Dõ��|�,�'^1�L f-?v7�W�b���l���1��ȥ֒���	N��:��\�9�ݭT�i.l-��^������:������uغlr"B3Pщm{8���6(��7�����:`4ZYC Ǎ�҂$�Ɲ -$���^�C�k��@i^�픱���|Z<�v��!�s�Б�̆$���y��Y�
f��'�
�Ru�Xz�A�j�O��O9H_(�@�
2��X�UǥE��l�>Vr�������%i��Lmrz\jˁ�%��(xp|�ƞEv[~A�(�t8R%����=�b ۽�����	m�T �9��(�)"��aZ\�>a	8M��0y�$[~��(nz�!���I6��ĕ�h�M�o?!V�(��?���Io�\�դ�|[���H�qK{",���T_6J���-�8;�@�=�ָw)<��	$�q�}t!�K�T{gg�R�0�,���f�T;L��׾\�]�+^	n���GK�U����}�m<|M3�+(�������Jm����C~Po��,{%[�9�A�5߱�!\iW�bEh=p^��R(wB�̄�*��J�̯1����T/�u�O:��)��J��x�H���k���4���CgηC�prϴ�U�<bҦ9�n��OB��}5�K�:(&N�Df����٤��lh�xVqY�v�T�~r��Vv������(�ߗ8���O�`���Ԡk�K���Ƭx�*3:F**��^�^p��'ݨ���\H�i�ˀ�Y.�H9
SVl��V�!��"I���9D�`f�i��˶h�\���jƮL.ϴ6O2�1K��3+��I>u˔O�i,����z��خt�� ^�L����C��[� m�SLL�d���r����SVNq����MX��Y9��(��7Ҋ��O��͸�Ē��j�����f����t ��vr.�̣+�_4-�:���űݫ}�V�U�J'>H�y��8��M�3�]�+����Ν��$
VV��]��]�4'¾��&�X��;��ԨY
���,%�l�P�1�V����r.:�/}���	�&��Q��N�^�����.2fq����l$�mx�^:�<���g�w�`��e��~���k�w�#Vom�'��ja+����k�����z�_���XwIбib���>G�p�c���5lX��D���;�X�h���%nT2+ᵌ!�B$�8�+$��q�ؕ�{��K�t�n�Ȅ).��
�����PzY`i1}:��i��
@�h��&%M�H�� D�K=�`�K}���|��*99E�������������m������#�G'ン��N���O+k?b'yrh^u��3����#h�3=pY�]�]<>���u}(M��b����fGO��\�V���2/o@�?Xus��Y��~u�aO��GL"�(~���^�E�!'�T̞f:����2+_�3|(�C	��������'DF�\7y)�07�?�7��Ó��3�&ۥ��7n��#�9\�3:T�����C��A�T>G�p�U�.[>sl��7 �R{�+]�w�T���m-�� ��P0��N�6Y�lkS�����2��:��|��+v)\�.����_`�nw��*}�n���h�	Z�J��tP���4 ?
�jf$e>�}��,M6���2O���v�c��8��a�N�I����L�"�B҉wU�0p.Fpq��3zǆ��K�ݷ�.�9�!e�T1J�]���x�&/��#F���K�)���V��VwO��pD ��,	���lB|���W�9a����F7B)�z�-�ڄ�.M���� ��)G�`6q\����r5���b`i���	�c�M��bS�H�Br�+��ɐ �M�����9�L�c ǧ��� ���O�@�3Jy
0o�#r��t�,=���ɲ�k�#}]���$�={�Kw����O�Ӌ����F�!N�>6&��q���ة���.-�ײ:����ڨ�ja߭?�1IX�U5��
�ȅ��s�Q�.C�
��i>n��k��$��
7AΊ�H{����8V�� ׮
"�綬
�� xЋzPc3��GL,�A'#���q8*P��ҫ�9���AY�?���a����Y>�´�@C|�7���R�ϒ����U-��L3W�)�;I�k�3�&3�II-�Oe�x@_�ZOPk��;��=���jly����P�G`����;/y���J~<J���9��m���Q�ySqb�sR�
�iv��I�z��4������E�K�a�Tܝs 8��.����nf2-GG�5f�. S�'��&w�ȧ3O���ɟ�k�o���9�ѵ�C�U\~ QdT�dĹ�"�J�
Vt��ZjƨW@�L�2��]�g��'��D�\a惆�~�5�8`����ĸ���G�s~�58�I)?W���+�\�Yz�Tdc�'OTʶj9�ퟻ~-w���\}��.�
1�pP����9�c�j:>��e��Q�Dk6��Q�����3O(J�RP,��!�3k5�Z��@��W��,�|�ħX�����d�4�e�e:x *$��Q�7T�rN��0ʉ	n���+7��.I��~���ږ{^�!'XL3���x�R"B���o��c��A�$.5?��ݹ��>���`w�����<�*p�@X�W'�D"������U�pZ ~��cRS���c���� ��%>�c:Q���Y�'�V��Ɯ�K8,����#�V��!	��ܐAZ�^��y�9�6^]=�Y�]�w�]�V���)�Q^���1 �	�"ێ��O�ȸ����ہO����@�h��� K`��`�⢃�����9�S�Ooa��Չћ��������:�����R>Ȓ&�>�&Gr-"������v�:��	��g�h��!� x�$3�������#M�ym�� ���5pV{.��H!m����V�噋���/$���	n>_�RبP׎p%~`6QT'mlM��w����s�֩\ch��dZ��M8�x����zҀ�.>S<;�΂�G�^q��	
Q.�[/�T������e��.V��Q�O�]�j���DK`p:�/�,z^ܘ�S��V��
�D�~H�����C���h�YMެ=&ƻZpG �3E_�)8����|���`��xp � �%�w"7z��X�dgWfs�^*M*�vE��� �8h�J�I�1�rh�\�wn`�w\G�l�� �;v�����óZ���n��q������
0��*�.���˳��ұ�����r0�Ŗ�=vHb5iڤv�HIl����ɉ��[�-�n^�7�ե��澢3�z�����	ί�5f�m���C.�/�Zi�.�w����p��̤��i���1��p��f9�YB���Y��`2�4Z)�Zw�$��~����(@=��S�Rd�f�g����ʿ��mE��Xk76����`B����֎����#�D��&�^���}/�ݖ^[�wE��Q���J�&*rǡC[��Э�C�u ����>0Ҹ��Y��jL��+�8��֦��H��H�%|y��Y��Qݨ�����/˃:L�k<�$Cf0�C8�	�A�C��J=����$I�V�Ӗ�kN���>B@�Z}.���\ cP5tl!u�ˊ�%�]I|s>�&�����?v+A�GI�K���_�<���g�ʒ��E���v @��J��}@O�@�5�A����d����Is��#�J�3S���uhAms�2��Q��H�Y��*�#�p��y67Q�!��/ c˙����o� �v]�7��}���וqK}��zX�H.�f��M�
��x
	?ܛ�F{���w=��'6��,F�PMƿL�z�1�DǤ��%e��g��/d���#�R㨶�4no�BM'P�r��W'I�!�f���.������D-����Q^4��j L��QCiRP�Ҷ���s��@��v`���/F�|^�����3��S(W~(�Y����8EL��)	V����x͹s̗��u W�� ��KůH���Ime�U�y��T�E�����@��N��� L�xdb�~;a��@$��/!qC}jz�㿿�Y�+���	�qQM:�]�xvܵ!I5 ��,gq�&�I}E� FI�̆Џ���ώԖLaHK���f��y,�P�7���;�L�J(P�8��Q|+rN�3TŢ�<�cf'IL���CF�G�))iU%��Ӂ5��2���d��|rS8T�f��ԑ\:a$�h(ā����|�7Z�j�vg˂*���.�� z��������ٍC���2�^�A��(8�lX��:E�0*~&ԤβK�:W�e>��ݘ��Y?��;�Z)��y�GA�S��G�U�
c��G���^�:!�J�s,�И�
Be�.+g��i	6���j�լ �&dO���5t2�X�'�����$���c	m<"����rls��t�o�EI�1�lL�F֓���@�-��!R�d����R�k���і�.c�AGra�U��2OJ�7��l�J���N��]J�����#T�Ib�C� �3h2صi��bl�����zQV�ݢfv����l�T'M8E��a�
�	��:M�h|n���ˎͦ������?H�گI�G� �{���Jv�M2E�0�����B-s%�\պT����]�g���
>О2��	;w��M�VG	�T!�eeK1��Ku��/b ����o�գ���-4�����/Z=����6L��Ѿ0��@Z|B۞��E0w�� '��e☄���"���8ҕOZyo�Jj�i�_�3�|;�ۖ�L��v._N~��^�Ҝ����ߝ�ڋn������k���?�0>���(����*ރg��TZD�GZ����,��>�M,��E�9M�����'{Mk��?� ���Q���E9����̵Y	�!#�ne� n��e>�F��S��`�.5Y�Dhb���Xy������c�S,�|Ɔ�-�����w��\��Q:��u����`^!aaA�/I���!���������V�y�u ��θ��PV9��">�R�L�b]�dG�y���~?���H؆9�a�fhvK|@o��V7	1L�L�����1�#4F��������M���Z-����BlK~z>�֞LSDΆ�k;��n�$��Y:�7֨�`K>�F��ݖ����;�"�C;��C )/?�~@�%g�Q@Ԗr�ʻ�=�Z,�E�`�j�@���Dm�E�׍��uN�=>���N�0f��������`;��"���������jR}���>�2d�� Z�"�~���R��:T�`�)1��l=wWQU�#g��0Yz��aɜ�����ҷ��9��ES^������!��EE��SC׿��VH�D�h`�/���7�m�l_[|l�!��etn�*F���A)�2��%ZWnR���혧;U�^��U��V��=-v���o�\mhc � ��%�U���jN����� �T���Z��3N����$D|g�X�V��h�#��w���@NQxgɖJ-_O۷�'r�[HĦO)cݱ`��d��K�� �(�a�	S���'�ܽ�8im�$��Q��L�hL!�C��������-�^�}td �ٜ��s-��0�X7�2����)��̍��^���8�>� �꯯�#��Y5ǉ����Ϗ�Q�i�}$N����(
��K�|�Ƴ�o����|��S}�E�ƅ����ДϏ}��������n{��zʕ1"�	gg1�|�P��_�e���pLi��I�RHOԖX^';���H�1(�ĕ�G���J]���)2�) ��pa��[X�/}�RE&���D���o�{Q�1�, ����ݸ����R�~N>�J�3tK��4�N�DP����(SV�j�F�C�%\���p�]��}�7C�U0[��g\���Z^
��谻��u�?}��x���ahzt��� R�T��H#[�JU�o���~��E�$�S�BPbl�ՙX�>K�M���z�����S���S8���R�zʨ��:[�:Щ�'�B��Wsج�)d{{�eFA� �2��ȱ���\Οai��9��8.��׳g�L� &�3��*�l=� ǳBc�/�`-�k2c�x�l�*��n44��k�̛�z�A�#�}�
���}�W��/&"����Ns���Y�+���/��LxI���CZA��0���!if��*E�j�x�b��'҈�D�m�����ƾRCڋ.�+��tUaI����w]^��G�3��U��S��Y[����J�Ы��`�c������=}dt�ط���JW���w?7���H�6���$LJ����L^�k�������B�ҿ��=��3?���?Z���Ţ\���u�	�2zM���_���`u�8mx��ۗ�������&66�[co sF�T�T�n>�Z����%;��1�+>P�7[�_s.V�� .4&!S����g�+q-��I�Ջ�^���l���B&S�WfX��	ԍ�Q�E�ʰ5�e�t	��+T���^5�����,ӎnϟN/�'����B1R�����v��3q$�Ir7��Ԑ#1}�@њW�-*0�n�s�5��I�^U�h��r�u��oM�䰽�/�/�7��������=���c@w��9u���Z̚������ZHJ�Y����<�F����o��jP�϶��܀���gm�u^~d�+�@ "s*�wHb�{`�YSF$��-_�J�Ƕ�xGG��}Fh���"p��Q	��	�bw�Ƴ�W`�y���!=
ze�����7R��w�=��|��#��P���'��1Y�x�^jI�bgn΢����;��Q$�8�W��k�ϗO�0DJ��f�bF*.Fś�-����Z��ߓ�JH�s��/��`+PiD�`!݁o���dF��E�6+�Aa��T�e��[(N:��:k"ʩ����l�������@hy1�_ ��A��o_7|X��)"&M;O��910Rȷ
�i�x��0���v7������Q��Ox����3�$I��ײ��xs!+e�B�d��0b���P���o���^��+|����g�^�?R��I'p�f&�ѕ�	�\���SԨ�]�Se%K����QU:oz!����1�L��ZC�}1��{&�n�o����p�R�*�H4m5�v�%Z�G=S��u�~�#��*zZ#�Ép�m������NӶn��]�r�:(;v� `b�Q��o���!աX�e~���\Eqt�i�wњ�zx�����ZH���,�2��D�=;UH�� ;ȅ�#ѿ��#&/�m=��w�K���>����O���ŭÎeB[�~ם�=tj�ğ.�0�_>�2II��������^PE��=�S,�T��2����96��:�M-!����-u ��Ц�mB�P!�N�2vt�L=9���\>s�F�ǵ>8��0���I4�&��c����3|�i����*Gn�����:��R��j<���1�٘��}3˂��1�RR���m0"d�rd�����^�LN4���<�e��Jc�;ŧp�ϛ��� R��`�%����Lߗ�<N����ٱ�f�����+���t�"^ ��\=�D�#W�5�ʄ���f����@�ω(��+T��z��˪_L��jH�����2.^��O/b�!�A�R�{ZiplIL����Àxٯ7Y���? �[����`S��������!��q7���)�0ɜǈ ���Cq���X�\��s�c_���-�k�.~�uÖn~!��q��|X����eG����]��~��{�д���=����B�Um� 4?m�m�;��Sa���2����]�-�o'��=��QP�]��k���c�p�����8?�
�͈��yU�*?㣊�"FFd�"�s���@J^0%��#�qQ��2O�V!v_+7��5R�7L"��[�Sj��	�V���,ʐ{g���j���;ź��\�p��*��� ���p��?�o��E}���&�� x΃�n�\������b3���r��~�ǽ����њ��B�;�0lz�����U��[�U��D:����6=oV m�'���]e/\��Wm�J��� ���Z�)�Z��W���!7�5`��-r7�3g�g7��g���;��rt��[)��C!Q'7NK����.��_�n��Zm�J��-�ٯڱ�y�Y�=��`7-��dÞFg2d��,�lŨ̷������It�ys�i�:�yUg3�;�dZ��J?�0���O7z�)�l�$�p#Θw#k��,�!��ObU���}�}��o��b�Pʴ3?w���5꺅|w�-���X�l�,vt�jn$g�V9����S�Ⴇ,A��b�4K���<�#��.�;F8A�x�rO\�m�岪ԇ�E9�0�_��h�<sC��7,��x'��L��
�Q�S��X��5�Y�6lؙ���f."̈́Y@��"�|ǂ�}C����=����W�>��/�����n�8R�uћ�2�H��H� ������e$�A�ӓ�b�{* �	�8=i�]�J���ށuу4�eA�+a	�Mo�"���G��jt|9\����N�Z�+�bHw֛�|���=�Qf�șg�3�d���[r?��8!����~�
mg�$�&�h j�u����=3|�]�Q�����h�F��f�5�Lo��c�f%H.>J�5��g`�|F�ql��z� ����j�゠��	��P#�ϻ!�^7�"˧�s� C�,
se�]���|����q�ւ��
�q�朽a���W�!�'�Ԑ~�'�dP��M&2$$1�gq������؇�<�t� ��0�����23]ڜ���D?�P3͚-��_�6R
[9�^DmHێ��{�C�H5�<�I/3�o�P=p"r$-�EU8�Lf��Ж$�bW3w�v�>~����߻�CS�ߵG,�תܙb]Ze��:�o<���K:�I;��?W�c �l%c)}�T��۰$(8�Z.�v��)�!	�/�����F9�<�����ց')�,&)��jֺ� e@�Q:�I�JF���%��///?7�̎]�/�,�UQg�E�|M���8w�1�r��'�D��C�������ye���[d5�"U���7fKA,�C�t�,|6�Q��n���5��t��3Q֐�F��4����X�%�c~�K���	�=��݈K'�y'vK��SR-���O�G�b�Oz鞿U'����������+;!C��5�;��Q�s��p�0�%����L(��C�-��;&�ҧ�,z���6�>A�͇?�����Z%��H+�t�jzC�h����0