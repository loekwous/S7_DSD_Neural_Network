��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w��3u�s5�]��B����k�\��"P ���V�f�b[-ςzehiY]��ĺ��n��k@�<���l��Ez���s�Ŭ�~1:��N�P�ӫ-�A��	�/P�r }��x"��#�I��j3r8���=5������ 2�� ��SB?����8���;dI��K��h'����@�X��ڷ�E��K��+�O9�x�"x#Uu�(C.�}ک�!�w�����r�G��wӲ7A�*BtԟF�;��1YX���g��&�;������7���ؘao�ꦡ~Z����"�YV���]z�����Y�1XWI���-���7˃�?��h�*/��a}��	>�>������1�N���b&��Q�V�k�?�Z�jL�$d:ړ$$U�{a����*���� *4`.�O2��Q��7��j���z�+����ɕ�N5��|O���j�O7϶�I����;��b�<����bf,4�{�H�k���~�k�	�� P�x8�W�!�o3��b\��^�Ǌ�gI&��&7|���Nܗ`�x�2���P2W�!�Xjౌ�BςwjM ���wDY1�>�?]ȑ�!J��Gw�e�Z��)���N\B��$�0�r�@3z"N�� }Ad�"5��9�[��'c&a!�y:^��G�&�E@�_� Ehƨ�hg��5G3{��������G�����	b��/��G\!ZL��	���|��8�F����^��)���5W���m��hb�Y��b-�Y���5y�=T�����92��D��{�4뗃zqs7�Lڡ�e�,y9ڑ�����F��$���22$Xo�~�;�*���;q�(+��	��j���bP���<�(��0�#L�K��E�iWW�H�(���\��Kf���!>�rT�·̓U�U���6�*��:2�blF�EU\U��h�kԔ��
�J�3'�{�b��oȿY&��,�>�S
�!�f��~K�v/�7H����UT��ꌑ���������`
 ���ȴC��KTqd���$��5�yj����zck�5�a�x�{���;:�<i�����B2`�w�/{�E���Ҹ+1ʡ����z�o�8����1v�4cdƜF�� ��d���e��b�y%� ��_8:� Y��:���p���=157��8r��«� 4� ms휖1�o;���~�'�3�%1�OT�s�v��N��@��y����<�?��j���ש�Q~t����S��è>߰�qԄ<*��5hc�+�d���69w���C��z�8�Hbn�*��?~�I���w5�O���(�������x-�����5+�	��ڴ{v���e�&���3̤���v|2�oq�Y7��zε�&J�4[���B��\a�/��[�#q���-���g�G���~/��f~��j�7[h�6���\�V8��)�?�h{ ���Z�%�ӎmY����%.�sd���F�^ ��GV5>��(�F���lh�T4)���e�.��\��[K��b�,ix߭ۚ]6d(ut3%�9b������B�u�x�P ��l:��u
�U��"\����rm�"�:?�Q�0A~!����X��[J�U-T��;N���>|v@�y3P�:1b(sJ�/u")�+�kJ͇X�ɣ^�5�[��Ph�%�D~����k1���p�<jV���yQ^���+�Bc\�Ҭ#L�U����NxmqlD]����WV9iz�OZt���R��׼neHc��ғ����o0�Nvc�M(3c��q�f��Ţ�{¢�I9J���ʼ�)4����9��x��Ϫm�X�@�������u��C8���ľNB甶��M�*�;3ieC8�)�Do�C�Osk7���?��Be�`S\�c}*k��xO��SL7��&/mX�eX#��&�|C���:���!\�`����� U1(�7�~�K�C��u�z�f��|j��n���M1"�A�U�~4w��b����S'AK���^�e��i#��5�]Rd�7@&�	��$��u04K��x#�JB��w�k�^J^WK^[Ȼ���,:��s⦩oXG��+�a-�׈�(���F�S�B�\��g@*!��YڳEpu�b�t(��.�`������Yb,�!Z�(d@���A]p*Z� ��kkO��9�#.�gw��D0��'�p�˯�WXG28��Ԭ�����M�}���2l��F� *pÐ��ƽO�iy�ˤ }фl���;K��Y�����gB�����d��1�'�%�r��|�G��6I��ڪ�\�G�np.�\�e�Q���NS�B�SM}4�d(��	a�%,H?{T�Y8Gw�;g��1�5��ĵ! ����9��4|9���^�^���tL<��@���`Ӟ��)��H-.d�k'U�wH����%o���b�S�F����[q����SOU����d�7���k�-�O�� ���[Wg:If�\2��6��C����>Fyb���=�%�dM�a1����J^��4֢��[+���=W�R���Ḅ/�V����s����Z9oA~�L藛�~z3܉�q�M��(E<���C$������Vl@�E���1�p�r�+?�n�>�����9`���8<����D�.�M�*R+��N�|�t.a'3��=-��g�b~�j)����g�R�4o�OX�u�E#YI_d��%�d�`62PG�Ce��zp&�`g�774g���րqE7P��%���)�]_���e��>7�B�ވ��>�=~)h��&Y��:R�����i�ق0��w��,���(���<j�nr��;��/%�����Z��^l���&�� +��Bdqu :��#ٯ<c&zRV2�Y�(𐽗�A��t��C�X��gzfp|ߛ,Hם�m=\��rf㴬j��:b�2A.X��[�D!��a�~�(��m���וgg��?op`�Z؍A+:5Qtřg�?��5=�����K��:��Y/5���1EFbm#$�q���;��8��7���ۛ��9���t��=���~^4�w?�U �ӊ޴����[�a��<A3P���^Мnͭ��5\�aS<j������ �\]2���c�gn�/V�����Kj�c�m%Ef�U%��߰&%�ǙfM����aY��܁HȄ�0��(�˜ � �H{��ni�H�f��Lt�]o����%�;ſR�z�/ j�!ʥ{��6�=�Ѭ]�\2�Bы/g���YW�:1)-�dS���!U�u�L�W>�#�_��s:ٓ^�+�*@�`B��PC�l�@b�ڏ�'�� i8���
�e|���; 2�H��#����3%�'xԭ�V��>]ꆹg�n�*���[)���ߌlH