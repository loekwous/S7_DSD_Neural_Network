��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�l�(���q�a��8`K�nz�w�V��� P�����"��l��p��2����}�iH��i�k��4'�����C�H-�%����c����ݮ�ƒ/L�o ��RD\���m#Ө���������tw��NA5b�7���ßS����2�+�X~듮K> �1p��M���%���|�8)�"���*q����E�x�-k��A��#����a 0�Ԗ~0Ghg�`,�i|v`����b���I���g �2|���KϦ�}U�+��t�qYBy"R�>D���tx܂�O3(�C�*U%f�[i��V�o���W�R�ѽ�	��Ǹ�L�8hG�]Ii��o�hk=t��zkC\V�P�0�{{M�^<	E�	��!G�I��E��/2T
�qd��HלgҚ������W�o/?Ґ���J|9�4��(:�zX	f���M_���j�)F���|�M+M+�D�j�eB=GF#�`FSF7�M��լ.|v��Ub��r[>?x��IOʕb�����5��X )�^k���q�����'̄�ThC|����Z�F)PjO�X�$4�G$sH~�u�c�p�������}y\V���Ծ!s�ċ��e7�p3)�c���H�V�,�+s����v��1$R�g���x��3	����tD���3E�[wI�P�t���5���#�8*`x�����=�m��e�)�B�gB�S\6��m��'<��#���bta2��[�9n gilZsk���8�S:SE��$P'j�������wM�X��]B�o[����j;^�&*�h��Hh��ł2=�#y����W�y�ʷ�Wd�7X�؋�KD�(gKJ�X�RS��{I��A�͏ЯoR���
�כa�p��G#nt{=���A	{b����m�p�^c=���Na�,�B��D��"��$��;���9y~4����nLܦT�G��'cُ6��8V�{������/3��x�۪���rZF�Fh?D��
U�z2�������M�X��P����_s���o�XE���)Ѳ��J`�����IA��1X=�d�)}5 ����ۅ	��ݣ8���8�]�(�ܿ�����t��XT�yxB�u�\N|�E���������:-�ݏVG�/EB����;�����\
�F)ۑ�v܄��8���/7�t#��q�h$��y�# !�E���ÓӞ:V��T�@j_8�|��n�վz���\U#V�N�5��D)�e	���Ch>�ͤ �'����13 �}���)�����$�����N�ꚽ���F�lv\�Z�\;�2��R7��s�s�urS��xwd���8;^}�9l(U�7�����st�I`5��6�g㗀��4��c
����Y�5�y���G�w��Lװڒ�t��̲(�ܷ�esX�{+pQCٝ9�V_z�)E}���{�{,�W����,�"//���p#�$�+���m�I�7wl�~�H��5*CQ�����;=�	w
`��UT�)r�i��W��8���@u�[h����~�%�c����j�
M[�����WA�@�����D�$�Kߟ=[L�w�Ԃ_�C�򍍧v�0\�E�/�/��E~Fy"�R���0=��ME��㼯M�}���)2p����B������L�42�J�9z}D��x<d	GJ|z��}�dU���A����'P�7ny�n�j�Sa��atF�zG-���Ā���!�w^\�7i�p�-�A��oM��y�A^�[�WE��񲚂-�~�%D�:{�Н��7�c���,��R2�7D�N۹G�r	��tm�>L�����W0�/A�Rc��R{m�Y�%g_Y��������*R�BP~��օ�mUT�Z��b��G�ɴ���-%�d����#1Wft���^^P��#�m�v��;�_��`e݈/�e߱���&>K�6�j��ko
&���ؑ5X���,���}D�$���hC���I�/5A� �l,:p��9C���!!��VS�g����8b�4B'�f�&ax���v�異��J� ��i�ݥ�o��t��ŏ�g�m�`��K�N����5v�i�Y4O�Ũ��Qe���H�j��c{��Gi�g G8g4�� ��\n�*$�*�e��v�n�"�b��\����K���m�0�=OC�	����Ϭ�d��`�۹�Ok{�%l��
	��cl��
FYB�P����\t'�������K^]HC�m��
PE�V盜o�t�{a�r��u�dS"��Zy�&!i�)i&k���䍻�T�
�z���fu�c5R��;��E�)rQPB��-�Y��u͇+|2]9a'��$�Ne��#�q�:%
��"��v7�2 8�roY�`�^$H&i�yBs�<k4��t��!F��]�X��އ9��7+Z���_��X#�6��9�RA�w��ᖬ�z3#�������j��\fjЍLi�U�GX9�n�V�	/�3{�QÓ�N����-6�A�O�_��ni��:�IO�D�'̝��Y�q<D��uW�#�C�\NJ�5+?iK^�
�=�ѩ+�2��e�%��_��/ǟ�EQj�km/�����az{�J�<��;d�&��K&\�;�
`���[b�K
�f�B�h�����W�[$a<X��ws�CIG`�ޞ<��Hfd�[�)"����ǌ�T�	)�����{2~��|7���Rs�u��&𶀆�/�3�Ӟ1Sw���_��L��u������G�S]?�Νe�SD6������.�tM=�E�)H���d�����J�`�_����H0f��x�ᰈ��BK
����ipIҒ��8Ks䁘���^&�8�
�K������7���2��v�k�6�8��\e��e�cN��xs�"��#�YPkc[��Z*�a��#��K5�w��nv8����s���E�,!�\9��:�c]VCMF��|s}5X�V�2�CE��.���D��!�|~�?�gq�3�ů (ɒ��_�e�څ�Å��6Y�����iwqV��%�3ĭ ����"ش`���a������g�2O������!A���o&Pz�����&��قI�Ok:!���/���=�6���Lb���-
���kO��������@>���Bz��7�n���Gp��X5��M�m�y;�u�ٟ��Y���C����g]��'�����}|�:����f��=��Fsƿ=��Y�E�Y��+	}&�A�}0/A��7��Pb�+b��8�:-Q�@rpV;R�t�-��DB@$j�r\YV%ZJH�ksTm��E-�e���Avp��"4�0\��(�[85΅��H��YS��f������|�Of��d$��ƒ&]OE$��#f�d7�L(�c%{gj\�V�8M<I��I��T����{O檌��g&�>�O���nLd3n$��`ar�܋�1��ݙr��,��QP��"�M�N+�ms�ҰA��;Zn6�6|T�����ܳ�0�Cvu�LV)X�1
^a�u��W��8��](i�֎˯S����sh��v ����=8�a��n�6�B��/~�^n	�i�|�ɔ�s+le����F��:ѧ7��Nd�w	C��E� O_y�k-hFq���}�@λ��R�܏�kv��Y&n�����y�6Dr҆gѮ�v\��ǎk�7<��G�P*�o�vy��lU���i�s����3�M�-������W�H�8���T�`�0P������G�u��y:=UZ�\��v���W��\�ǃˈ4����ǭ��9�%�`�U�����偓�JJ�~�Ɵ'��U.�(\�L � �˗h��{�jBv=���q���l<re�(�� N܎l�y �^�A�]�����]}\NE�2�AeZD����n���h�;>�{lMj�y��ߖ������Vpd���,��;@ *q*�jz��ɞM��f�4��o��O⭍sK���kYL%#�G&�	ʅ�v�ϙ]�L�~��w�g��4y,\ki��$"8>�ɡ2�+�8�"���y`�R���Krtc� �X��} ��`���S�(1��KZ�l�K�/���U���) ����}�d۱������۱n54!vN�,��N3��~N�fE,���z#�`�s�{u�R��^�`�U���꽍�;�{KM$?|�L����?��ýy^{�_c�C�SgR��C%�y�c�$\P�~��ʉӹ�����V��r�����K:��[7���̂�5�f�$npX+�#��i29>\ӓN��ld"?I���%9�u>9�<�6�$'�<��׻V�	=�nE��8W���V�_�>נ"
���n&���Wn\`_�#�j_!�H#Ն0����z��?�^���¢��ې�OL���z�lz��g�A�+	��y��NV�&sS�M��2�`g��7�����!ph��i��Ԙ�����e��x|�e�B�@y/dP�F��*`^�fУ/�m�G�[�5?�mG���4�mxC!$6��p�K<	NrS|�mM�޽$�hh����/���dVQx��p���D�,\D��ݜ�ꃶ|X]c����[������jKZy��/S!���9u�	���ﱲ�tTiB���P6�U����pA� �>��Oa�kE�4C7���
W�h3��[��y�+���5Hb�����OhaɭC~��$��[��'�0e�T�v��1��,y���v���‿�^�D��e���:4�8jA�2,cВ����vHeb%�.�A����r^I����z�|@���_���H~����M�2xo��Ho�`B�0��8d�e��J��h�;�/��x�78U�����X�ǫ����E�(@��3<p2��_\�^���ɇ �����;����������æ��|�آ���Kr�x�'w��� �Jg�44io�4)�<�����n����$����${�ˏS���yd**�ehޥ�����}%*�.�A���l�#��e�Ǹ��F��pA`�,=��yz>�A
��D����f �{�~�|�b�/2����.��>����Xy�7�nb���"��4�j��\4H��4�yr�<n}����JJ�ceC�wr�U�t;/��9�_>��Ƕ��H"
*){�En�^�KY�x�ˈ
�`��t+�YN���q��jY%���wdI���D�S3��L��4p�+K4�:�ߤ�ҩ��0{|���	���ŕ=js/��u�MI�s���W���%$�!���t"6�s�n���L�m��k�@���
%�'���d�*>8�~cco��.Śt%q��;'e�z��;	~��.���� �Y�,��ss_���k�/�4W$R2b_�dm@�b[>��	^v� �&��@���x�G��u��'��FtJ�K��O���%�W.�޳$���!.��"cu$|��L�X��h�p�Z���,��<�r��˽��#�E|Rv� ��/�X��,��w��|��Nda� �*\�}Ūr��?� r�'V���E��2(��!w.�l'����N�-=&�ӛ�݅G������|���N������z����,ټ��dʀiR�K�j�{F��g���%��5[4'�?����Lj/����~a�4�k����?��I4j*� Н���-r�z���EwJ�)#�"�����Ñae3���@7�����;{J�3?�gIU�ᒙ ��^�g����n;�>sX3�o��^f�����F%z����(@�Û&K��o�)=���S8�WHb40f3l?�S	>����_@�1��H]$+H�H.�3N��6 ��
n��u�d��~%͹��e��a�{�`���m��/��iN��M��I�X�VR4�R��:�S�8n_K��40E�9���b�EO���N���5�(���t�T�tވƳ��(/@��oW��n��g�mDb��L�t�k���ϰh��D��$����Z��u��k�4/�͵�KM6�{�4i	٨���x��X;���M�%��ޕ�m�	,�S/ ������m�u�5x�E_��L9����4f�`͛������,n`�?�ĕ���5�iwXM5�me���=ua����:1�(U�XB	���QA�������5|�Qn� ��U���*�d�<阦�Օ�+ m���3��4v�&m*X-"$i��O��hAȤ*��fِ�}Ie��~� �i��SC;����x  �֬�.YO�3����Z5-K��PKL�ڵ��f�����U��`�}���Q�׌����v��J�\�T��!��t�/�cL��ҁ�CD���n��qp�@����;J�Ɩ�㶃�|��-��@a�i�iQy�Bdz�J�R�0�J�f
�Y��0>���4��{���r��@����uW#�(��E�!�m*�u:���^&��L�y
R)��i�XG�`Xt���ڇL��ˈ���U���c�������Id����dG�݊���8L}���l�rf�
)�+P��������IK�#��#qx����ӣ�qj);$�t�|��k�7G�i��͟(�zq��'��ʿ� �{���ur�s������D}B1jO��zZ>gyJ����;F羣�p������ k�U�kq�%�20[^n8��r� �ݕ*~c�*�L�V��P�!��*$�Y]
褞�l��Lrl�@�v��t�� �?�*vu�_�k1���is�Ҕ�Ł�gc�3� ��}�:;��6�!���J��PeP�6���%��Y���o�υTڃGaJ=�Hd�"��q����4�eH��r��tT�- m�ևL�'�J���a"��%'`��F�����q�m`Iduh�Сy �	n�]�0-?�0��&��!G�����n��J�:��w@���{��烖�z�}O����7�|�z���]��! ��N��d[Y)�~�#aUDe�{94P��$/��D��Ҥ9��0y�������G���t[ڹ����6����� �������9��Z��!c��#33v:�A[�º�j��K1�p/ U������v�8ֆ��%h��}�ʗp���̲����6Pr�R��Q���|����{m����
�t���p0p�EL/������K