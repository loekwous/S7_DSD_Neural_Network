��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�=D>�ͺ����v_Ȣ��n}���-�mp[�=���'bf"j'1��Ӛ�:�&_�x<-61	!ma�]Exz��l/}����!ֱy�г'��S�?r��_}.��gM�f���E��Y�Dݔ�����~��A#j��QRCIP̚X���u��)��� �H U�8o�.���P"Y����bh��RA5P�w��ޕ���``O%��D�d��]h�ܬag�����(���|���|ܺ�