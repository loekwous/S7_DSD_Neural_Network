��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w�6V�%{��xb@Z	3���ĥ������2�fU�0�;�=݆�>,}��	�i�����B%��q	%���8n����o�k}�ť�7��l��� ��}�y�0��4�M"�!��1�p<v&X�=9��s�BP�眷��+�u�����묩�&��i���򥉿/W�V7	�*�@��y��ɀ`w��'0��M����DlM����U���et7.��jj?V��{��{�ј���랢��m�d�Zc1�)����Nޏ�}xӹ8QX������i�->��N���|?cF���Iz>8���_v��xki���I!�a�������H���;�aa�R�M�1rS�Ak/��sr&!��;���ﬅ�t#����o�;�eOO4��]�?�L���^��h�<�R��ښ�*�<i�$���^#�V�c�G� ��?Rt���8��A�f;&#�u���
�u�)}� ab�������bȸ�"^���R�2!9iQ|�C`��P��*����-�~�Doj���20p����L�q�����t�LV�/����]X�0���]�AG%�[����\`���)�yG`�Q��E�X��6L�?/B� K�U�Ȩ�/�7!CpX��l�)u:yXeGm�/-�$*Q��Ȧ��k�|�v0���1�f���|j ���?>�/�aew�%�KO!�:H��P%�²Ǝ]�-�#Z�%�O ��!w�r��Y��P�6��?LR+Ur5i߂l�>r����-2D%jκ/tY���K�St���2�����W�.��%�{Ո/�ӛ�[4�I�"X�;N����2<�3Ymǿ�C����u���j��yB�}V{&T�7�ْip�:'�\q��`&����̾$S����/%�x/��c	K�鵒����m���]���|�Gsy���Rj&���$\�g����9� ��pg��tR���(1�2{Y:b���؟��8*�휙�p��Ǔ��Q.�����K\kLy�d��J�k�ț�sƢ�"�9%Z��(��'����;�	�캮�5�v�C������
qz��a\�HwziI���{Jr@�,BEE�(ڏ����҂Oɳk����p�55����w�w�2�9x2��Ê�'�E	8�huw��?H��2���\�\��
����"�� *�F碿BHI+�K}*���ׅ�h��u��ՅHD �/��vR��h�i���b��=�̝��~�"�-#�G�1�FZL0M_uMS~Vk!8���5/ֈ���w*v�n��%7� �����=	�}�Kl�ھ@�sx90ַ�[���ʅ�;cԵ �ܙ$?�II9���e@��B���2���"��+�������̣Q�6?�V�G)�C��GG�����g����|���=�IǴ�Jt�D��̬ʨ:���\�K���}z�pAz��b�M��!��Z<�h_�w���^WX3����s��.����dv]��8��͘�v<���Q�R�7���Sf��Bܾ]��.B������u�!W�眇>1�����:�2���$*5��`�=w\�we A7)�p�!Z�2@���l��\�;�51�͌?��Ҍ"�s�&C��H�g��.���"tb��T��B��]��1b$G��$����(���O�"��&��郵@MN�з$B�8� ��go�s=����/7��xu��Y��N!�8���
����5}_?�=;њ��g�ǄT (�>}�:����l��&�V�W�2qt8t��if/V��"|wr��6���E�KC�OFLÎ.(?�5���{ތ
�K��������$<|�J�b�������~����E�*�L��L$�w��Jgݼ`Pl���$�[Xw��;G.����Х���Ơ��AJ����U���a���I��h�~�EZO��WZI��h�xq�E~g:_y�=3g��|���r�Y�ZF������/�Q�kZ{"I��b��8`+4���̷�)�� q����|\M2��M%��rC��c_�N;*\�2!k-����h�+�CЦ](���+"xXn_�q���
���r����p����3d:��W��p�%��r�;���K$UpS�+�VM�M�
��g�~� �)�s�<-Ƶ�B�L���:��s��;ͥ�Dh��.�@%c�xZ��=R�Q����U"���ʺ��}�W��[X�
f��MAN ��y�=�y�e��u<���DN�?��6�n���=�T#צ���.-JYBA��^�_�,R��l�BzҘ�HP��!>KS&^օ��������q�1�8�����i�����H�B����W���u�����M�z��7��8b���=�|�����ȝ��i����������K^t�(��֣j��@g���-f*v'����\�����o3^���4�[� �<M�~&��r����N�I�1��rP���� �VJzN�*����� �uz��!JR���?7sd,�������!��꩏��h��E�~swY�`�[�=p�[��4���/��@��Yk��A�F,�'ڭ��l�;S�����f�V�����q���(��"r5���n\������K�0��� SF��\T�l[	,qX����� auk��GU9$�c�x�J`[L���e�\Sю-3���o0�t���5F{�.�Zg�SL �J$e���9�����H��E����!Ǚs�4:ޏ�%�����O�z�+Z_$�1W
��������h�p�dD�u��*
~�Akp���!�����$�jp>�̧����SP��?�k�-0�JL�T�0\����/0�G}�Ƌ�Q�|�9�rw�4��]즍�E$�P���I��9��E��?�kb 
��&��f�`oaRh:M�Dj�����{�Ixꮭ$�\����H�+�<�i����9釕a��뾉}�������N@�ba��;r�i|dS��,˒���F�pB����2<rܺ��9�YҺ\*�|0J�����a���aδ�F��^DO�7���_l�?û)��~�Z޹ߋ껨oa��x�Fq{v�_5�����^�]��9����g5��V�Z�5�}�y��
��'}/��\�Q9�ԗ�!МT���#ݫs�QA?�J�'��w�A����]j��RM�ܗ��u��OO��xd��^�.�����0 �g�ekE��!����GlPEeq	��ŌY(�1x� �e"܋$ yj8�P�a�##���$�^���֜�Wǥ�4t�q�f[^��\��&�w��������U�}��XvC=M�n�y�i,��te�c���<��6�{+?�:�BWP���r�qrEE�x{Q0]GG�A�J�L˂@���Ǟ�9���F5�Gve�]���H4�c��\����=m.��v��i��I�;:�2.�E~�
������NiRaD��d�4���g#!�����u{(����L��C��W�]$h�lMn�\M��H�D�|�oU
}�k:���P��rJl��W1QP��o�p�~*�bm��rO��+W�,^��ԕ�Y��\}��{�c�}���_���-u�檘�Zq�)!�h�7�u��o����p�а�a�ފ�X��d<�g2؉c���0A��@I��'�����p�B���)�AWJ>��������F)?�;E ��wp�����(oHl��Ljf��ѼR��b7�B
�;q�jB|DW��aK�W��#���촵E�M}��pR?�H	�Z���"��q�2R��X�_8�snY�����g��j�o�y5�k<,���Z�,[G��E�6� ��h\��yT���k,�����d�Zj�}�A�m!e���ҥ��C��>u�8!2�bTE��'we�NZ¥�o�rq���]jU@u��� 蚱���9<�)���z`gZ�\.��-30�O�'
�!��,���顲5>�X�΅a׊w��	X���܅�{D��yZ԰��aF�T�D�vuj=�B���.����R�.QE�=(c������ܟ�Lcd|�­9Ϳ��1{�RGRG�|P�k���EZ�����k�Չe�q�*��`S$�x���O�BV��Z��R�f.�,��� )����P]I檛�C��ح�$�f��DUNZ��灡Y��u��
S�����!X�9���^�@� ����Ы�I<��*��9�Q�١��$�ns�YM��iO�G����+.v��gg]È2^�L��=���7�!�*���Ӡ������gT�m�$`��S3�M-��}8���� HƠ�^�)е���N�����-�������Tvq���8AG�rԧ���:Zŀ�&��D�Ns��\�"l&��������hݓ���1�+�m���S�UH��LE���?M�񹬻�޳1���ww�ǒS���i�3S��2�!f��\�x.����]��P6����׎��g�����F��	��u�?�j�O��g��ތ�&�$hk$N�f���u�$��� ���-�	ü���;㓘kW�p���2�f�:`ω8x��D�KZ���-�>;�'<�q$�x�1,<	=�@GIR[ak���jo���U���G`�YҺ�)��ݖ��i�ǲ�e`4]����D!��/��{�K��\ٷÍ3n	�b�ΥFXRp�8tӾsC�ä��^ю�CI����%��j�%���P#\l��'m�!n�^l�e�c��.Sj�Ti�f-�1Z::L�d��A��\��*D6��ɯ��B��iP�������{]v{�(D����#�;�יzs�=�}N�~��h~´��A#���>6��O*KԻ��["YФ���rG��}�@_���rqc�9.��y�F(�O��1����R�!q�� .���.�-��u�����%z�I H�"x�)�Y/F�6�V�Z�jNJ��3.v�=���u >N$��aJ��n�o�A;����O�]��~�g�B�x�5�0��i��IB�3JA9T����~��`�0��>Tn��xX&����j���*���k�
��9�$� m�5����ěa �7cc80#��1f;��� �����=��
�ƃ�=Qfv�%t����XL�ɩ�\	|���2:o$k���?~��6%�	���-��Q�~�?b��[9�L�u3�</s��V!�'�8�HmB���?]?	|�(�^�Om��@�R�2b�o��^$([n�x�ʑ�.ȑ.����%Q�h�v�=&S�T #�Nh��1�%l��v��M����F��r,���e^���bd��ƍ6���l��׮�2#+P�k�^��$�&�u����hg�2lhp��j��N/�͛+�ʮMm����X��H�,��ޖ��̴�T�s4P3����u��!mw�	Q^ 
�Oh����.�[�����+�`6-��,IwE��S��?��l��A�iK����b6"ae1��,�@q�&/xQ��[�Qx��MV'�qy�}�K�k�Q�*	�Ǹ�4��7��n3�5z�;�d3)%ݣp����]�XQ�U�7�#�eV�����.R�t�OV�?� ��@�C��hgc�G�����:}mǍ�ž���G̝��㮶�3'�u5=�B� �IuWA:�Sߨ�=K��/|����D�6��i�\�*�*m���Af��S�p�0d,�r�t{pE�O�s���bc���D�5�SKS����x���iܯ\B������������bI���a�P-��N q�=��ҿ�]�Y�d��w��تBy��ֈ�<68$-)��\Ǡ�ޤ��A��b�;8�$�GxR<um�_n&p��πe;�#~Ybr8V�Ya�v��@���ߟ��mUR�,��"��y#�������Kc%�B������z7G���s����p)֭M��\���&X���qQL�kO��G�?~q�e�A�4\w��^��cb��.�e'��� }�:�e	�UF�[K���|mJt �u��7��\�dc�1����:� �=�0/)S�L����c�w4�F�b� �S]Dv�Qz&�^]�;C�x@GF �4�z�>U����]�I�|iz���M�V��>q�()f�x!�*�:s��b{�c���L[�� &6�N{A9��'c%���P�G���K�VԤ��҄����J�Ny"�|�k˔����a{�1X&B<�6�r�$��c��R����^O/2��ׯ�B��w� �)��M`KN�b%6�(�Lߨ�#$�c��=�ϩ��`�����r�ͯ��qM�MQ]6��&���ɹՒ��0FKL���E�>�5N�ܨ��y�y����z�u��c�Q:?GJ������_)���]I!���'����3i�	L��_��u�_�� ���d�����U3���CJ�\9�jp~���3nQ]=���=��&c�>m���rA�9��C��@��ד:�JA;�Eۏ�Wk�.Kw�JY����C��������|K;tq�ر��q̚ QD6־����"?����n�����;���HW���D�.�ƙ�07B>�=��F�8�3nt���B��j�Wϵ2<�+tZӅ�|�آ7t:O�F��
�w�����B%��V�)+��"5�p'��	Lq��y��.�Z��a~�"��{tb��w��^s���u�����9S.5��5���ۮ$]�ɇ0$���.��]�̎B?���Xci�{�`�>�����J{��|��ۇ(��#�kM?k�|'����I�sSYƯuz�-'|3�i����� ���&�US�fH� �_}�����4�<@VR:6V�dv�?��Sn�C��E!I�*|hT7\����dd�h���tho��YL�߲���7Ǽ����)ݹ��H_M����@m�_sD":?~F��>�6��[���6�^��f�j�1�}��g����T�$	�����"����t��\<�ӻ�BG�}�Ƃ�LBF��u�q���t4T�|S^�������7��[,�w� �­F_�Kn��ם�U I0�L�㰨�8���A'�� }�Fn����q�[1��wZfM~re�ui1X�M�O�{�)��lo�8�B�>����s��5�J���n����xw���*�hgޘD�=�G��o9�����p�y�$��Ȕ���/λ$��GU� ���"��qy
Z����I��¶�r'�h:(�4>��r���;��rv#_,�ݚ�1-&
�G�̴��z�u;o�I��^���%K-o�$v���]���k��!O�y�p�$��	���_��VT:����j�����.�f$^�����s}+�$�O��E@��m��N�ǎ������M��t��}{��-u�~Y�(���A�BH�ޞ�^�F�����%bXt�8�ʯ,�*j��5-%�N�|��T=�ػ������&����Y��G l-i�@WVn�+%�D�$���+��q�H�w�H���}II��5��`�&#:+���}l����yjs�40���u�J
����O��.R�t��m'�abD�YD/Y�D��pS�{\}'�0ʵIL�<}����: ��%H����H/��n��(�7,
 52���iB",�s�K�o����8V�K+���(+�/J�����%������Q���XU�D�f�	W��3�>+Ac��\�ͣ/��A�	'�3i�F��$|��w_"HcT$�`��Y=��ž�����ܝzGN�xG�B&˗�c'#��4ݔgZ��ۿs�L�Rk�ԾG�	[+2#}�|왛���4LX(���]6�*b����_���qnp�8)���<I���x��_���u��߈P���S��4�io=�@���Fb͞�j:�a�+�̝w��al��6����y�b�)9��X��WHH�|�L���7E* ���gTH Y�p1��C�Z=�f��=񭬂=4�9�
k=���g1np�h�h"���yqץ�?-e�����7B�)W�K1��_�V�l������Rٲ921�5�5���)߂2^���\��a�k����%������b������y�IHX��F�M�4k�4Y'O�D�}<WK����Ls�����ɪEUtpύ*��3N;*�z��`(1s@e��Bu�Tr��>7%�%BW���b�P`�1w�h�h*�ȅ� ҥ�	3t�*:��:B��R�Yx���)Y�1�.�L;L�Wc��Ï�B��*�bl�q����9�������]�H{�@ڿ@D�P�����H��������ی�����T꺃R=1H������Ӭ��1���Oj����0A�]u�a���%���ˡZ�X�d񵎇`��n~�2�X8�H��h��x�.�,}/V�A8�co�2_�"i&������Ԃ0s�qg�D/ � ~�>#[ʺ=��'[���֌�����)�?��3�i%5�kJ!����oe?e��!���(�D�!v���#�R��H�ih J_�Jdߎ�Xi�l}N�Љ)�W�17:]��؜��V�Ԏ�yI ��!͎w��o8���N��T/8K�lS=�(n�3��ܢ�O����3�M��KrE��#|��9|���9�O~�i6!�ά2H�i���7ѣ��F�^��&�4�����[|�T/Oo�"�����+-�I0��7�I1N.�R��S�x^����,oA��aNN��[�O�r�C���Y�C��nbP!�݄�:�sp�Cư�/cU}�L���G_�ښ�f�/d`�졜w5�k���@���~�Y+�{��:����9>�F齵�9��C˿������<%��Df{�)����-��-B7�D�1�*q���)�(![z2G�a(|�4��O���W̶N��f���sn�7Gb� �$+f�B��g�S�
J)fr��>%��4��5�/5�*�]�l1Dp��K��ezɏ�P�f�� '�4�à��	���W�&I/�W������]ͷ��(�:(���Y�sE>>�0��}�m,�}��s�_{wT4	/�c|�w�JG�E�M6־Tc�L'���ﬡ'�C#v��,�a��#�f�:%d����g=�vַ̀m�<
ڔt�d�R�Cłq1�|�s�8�$~�p��/9�d�99�~�D>�.���pZX�G[����ѹ���7�B���J]�y��[.?�"Sq4�((�wU^4��Δ�U���(t[3�U]�A(��(�܄��<��#�:�Q����w=�Z��N��+τ��%G����C�\��F�jz��NGo��q�ݑ�4D�P�0E��v�zU���'�ݻ�fh��Ei�SSM�f�硊6�ܺ���ϵc4�Ƚ� u��.���l�x�ͨ��D�!� LL��C�?Ps{k`�i#RMr�?"���ٖ��`6.�$�gV|��'>��2�Q�B؆�>W|�&ѐ��n��r�����O�u�+���ɏ��#B+�h��Ï���U�-}��� �!�9�ƈu���+k�𩘣��V��2�
3+�f�:W7&� ��J0I�@K��[��UQ�F�#:b�t1LN�M��PY��	n�M��1���Ќ����:A�XD�`&��t�k��
�ک���km�]�{��P��%/��'�`7f1 �br���ˏx!`j���N$�;I���:�-^��:�U����ԽC��X����+E��:.7d4X��[�".=��OA˔+������V���z��@1�<~���rμ�h��&������sT���������BQ��$B�!�fn�k�F*���r-���]��V �����;5�����2�
s�ͦrc�3�K@�}a�Z<��	��
�8�w!��T�Ih�qk��l8U�@������彪�J?�R15%�K6��u����a�]J^*\߷����!���������w��Ҽ��R(�ε;��	CB(�M0W�r�ę�Pf{75k����$5���Ǉ񔗗4���1��x�g'״W����Z@k��	�A�om����C/v6�z`��V�*8
���sE'������k�/MaI��o���v	���6"���f-U�7V�!�DJ���&�@=�����^�CgJ����{Kb��+{����ԯ��HyV�>,�K��~�P}m��O8�|Ā��� @,�`U���}�O��U�ڵ��`P��UG��3�1�&�UO:��	P��u+g�۶a��2Zz M��FPy�����X9>�j�{��<�q�ψZ�J�%@"�%�.FD`*�?[D�RO���Ep�%>_��b�i��O7s�5�f7�6���ډ�E7��(��!H2��v��G�B��\���u��P-�mߺ��%F����Lư�S�8O��)�V�p0;G�Պ�ˏ�'g�M���o��	��Å����ݹ��P�j��4���Ů2�������$♨I���{�l1ŀػ&e'�8����A�����4z�R����:��U��Űᓏ�]��H=��n:C�����8m�W�<������Ґ��"RH�5�)� ^���8g������Xd�-ޣ�qRxZ�2'���%*le�H!+[$BmQ�+*�y���g��C43Np�[��MS�I4N�T�w"g��)ͺ�ظVN� �F7�8)���h�[���x�V�>nu�.��`2��>Iچ�G9�u��h�a&��[u�笓��|�P���rŹ����Q'�9�B�(�"1en�6���1!�][�<4LKè��HO���_�9S$k�15�Q��0��࣢�V�оG)J�a����ٙ8+|yeL<��t���j�7�8�P�u.����<��j�]ik�`�ڗ"����ܞ�pv�QBJ��4-�q��z�҆M1�Sƨ7��o� �~�[ipNA%߇�R@���VF�
=ײ�葉������S0��GE��ۢ
�s�:��Ǐc�n ���{�̥�q���Uo�X�����զ��E�lN�N�@���>���m��+w(�!HR��b�=��q8�$}Z����;����l�Ǻ�oֹ{����ǟٓ�KN8eM�E���V��;����2���vM��*te���������؊�T^�(�v�s�(���=�B�ʹ�t(��caIz��
c��錹������M��Aʇp��䫠�Ɓ�ɭ�O=ԁ[8����ׁ�r� �����o}����$��5��"���*�{�� 8��e�pȐҿ�n �����#�d��~��{ʳN�u]o`3�'�o~�8m*^��?�����Dj�A`��i�%����M��e����/'�i^����$���^!��1KWgʹ�_}�ͼ�u���7�,��u�9\̧�s�uj���2U%�0"#M��c�{hCM̢��(�Y��&3V�,����جמ|ִ�NjOW�j�fv����/K�2�����@�4��u��F���jt�'���>��̒��V��?9rm�v�g�V�·�׺�I�U�GxC'�`=�,����~H1M�^�J(E��;Ee1�k�����_�e"0n�zǆ��1JPI<eY.ƞ�CQ�ɯ4���y-����4�d�;��/��/N=p��OR�;�Z�T��8�y�U�4Z����ذM~j�����c���i}��֥�$�x�C(Rq�	�&���T�Y8	,��M�WϾ���
Xe�W?�
�����|	>����'uH@�G'#�s����k��5w�۫�R6�}�@|'-вi/�D���@�t�K�r-���s=�X	o�����b��C;����+v�3.���	�-۳�m	
)G��?�Vچ1�����x�ȣ�X��b)u�4  �*��}͡G}G�Qf��Y�I<��"(;.�H�(@� �&�(��W��h�T��qa��Կ�y!595}��[N�oB�lV�K����L����K]��F<��I�ȍ�c����Q���1�)���+�N�]0���HqB��y6���2�^�0�AC�
Ӄ�p�m-e��x*t�ԼP����K� ��q�j�лa��}X��3���B�=~�8����A%����
���.v��]��� �d4�����IX���?�ڧ<�j�^���a<�-l�o�n󰳚c��&�7���ny�,�:�0]Ŏ r�6B�	�G{L�*�l��n�Dm&%Y�~���aO��/��Ǣ|P�w���G�=���k�ױ����wP࣮��k�U��%_^���_�G �Eҿ�! ��hs��4Ʀ�H(,�Dk�0왣&6�gE���}��i���B�<�;���k�-/CI}�=g��u@ԫ�q(��U�37��#��.��cE�A`���}]��D�!&��$�+�ȕ�&���5��3싈��6ua��xFk�]t���;y}�Nd��b���!�y="IcHY����u��u����g��D����R��`��Ń�X�B�ɺk��.Bl�+9���e��?TG�����Zp8]��M�D}	7�:���9�ҳ3�"���_����UU0su��:�|��:�h]NW}+�����v)���m��	S�P۠��ǥ�cϝ��)������r݄00�A�2|8~!�-3���D�(:EQ���o`38�¯SyyO���D���ɾ���Q�r��^9�e`��gq�1n�3��U�R�K�cI��K�bU�4n��q��0=xg%N�ĥf��w�n��6kV8J=�I5��Eg�t~��ѝ��m��ٸ5_�+�D������u�\���<N�d��C�_/Nͦ�Lb���Md����#a�ϼr������}L(��4%��iR���"��F��5u\ϛ�M�cw����a���]�MZW�Z�o�ؽĲ]�e���V*��G?���;�.6��3����Q,�߸;����qSӤz��؃��M��5��m	8�����r<�d���ε>����W�ct�[vJߐ^D��|��^]�ڲ���aGM�����
���w��"OX�5����R|0#)��P���5� d�y�a��UTĬ7l(a%6�T�j������Ȅ*ǵ(I��t&fW9���&{X��n���H��5�m�6U#�MyQ��9�]���	Lݾ��F�"ܠ�����b麎�Z��x���at�����f��R��T����hx��
�-�7�(���_����Tm�'���>��[*�o�3�zn	R71�ܚPp�+ŖH.~���.��x@��1�zƬ��~N�x̲�2�B�o��\����ѐ<��A��Ba>8� �E�x�dpn��j����(����=��6e�.���)�PtWo�mT�9qe�<<�|$Ժ��ք�E=���I�Ss��&�ep`������_���T���@M���Z~��?%�3��u�T��/���F�{�X\�%�y[�u}�$o���}&����|��4֋`�?��43��DdDB²C��e�jtp8<�$ٿ˨�&θ��ť���s[�n��ɂo�܁&)�zZ�������$�U �k��!�� e��*Pę3`0�Ĳ�3��;�rp�n݆,EI=�:l�Y�����U�H�`!�)K�i�D3�N+�ۑ���!(`u�dj�n�NIuҠ<;����ʞ)P�ɨ��b�K���KKZIe����,3�Ո_�e���#�Õ<u���g*`��@��G���͙�9H�N%���v�^Q` =\��)3B��
GXX�&<\�Ϣ������*JL]� �ZG�m6a��4s��`��b������&���-�D�d��u��}
���bm�h��\�?[t�Rt�L|�����-���m�W�w�nA���Km����s��	&�js�?w�fD�$ʻ���h��!Ԏb�	J5�%�W���A�g�	"��X��S��H�	�;�حPY	p�bP2�	�B`כ{8�۩˾օt.@����ҿA�҈tlUw�a�D\z���;�%�El:~tK�O�)YB�Fg��l菪���B�\��qY��Tۛ���Q��|*-]�R�1���@��cd�2�H��n��&��񂔩=[ƌ|�4�:W��%���9��\&�";P�p��/�����>>���+��7�4�p"#]F��ե�Ѐ�B��>q���wTP��q�4�٫T ُ�ő��A���Θ/$�g�K�C`��X׶<��b�����nw.F�xmW#�\~�bF �q�fH����5�]W�*��1�?c�UrEf8 i��w��8�F#�����@a�S<mxd�"�e��p`�|)קk9����R��
wE9}�_��d�in����a�/���b�nV�HO��~�)T4��苏U�f|�1�!�)���R��0�T}xN�7�:��^���O�ҺT9�%&|��;)��La^1K(m��N�Vg�o��<�n�?�g�-kKByV?�9�&�n �j�wo�8i������2I;������e����0�$���8�4ܳ�.���/H]j�������
�J�^ݘ�P$L N3�t.
�hX�����f�^ڛ)�Ͽ���[��i�G���J����q���:a|����?�4�t�2Y�U��^dq�=��^�l2�#2�8kQ�F��8t�j�o���Q��n���?U-���,2�*��x*m�'�h��`�$�E�-?��[�T]��Wۺ~�ۍ
�C; j�����vv�͢��4r��U�m�6Q.���xzI�ٝ~�]]\�b�0��b�����r�M��r�ߧF̡�	�p�]��) �d�=�D�+6G�s�cC�|J��1�La��|<L����ր`�z��x���Id� -~�	D����[��7Qh��-�j��*v�S.���p��u ��.���fH^�$�z�7J���C3ⴌ�#�=�S۠�&"�t�i}�;f1�^��N��d�sm/�%����qu����SrWhy����,�[@!/ :�p'��M�c�St�U��g�7��d�-\�9طf�����7���/h'|IO���*��9\Z��}��w�RK�@eW�󃍴q:S��n��TE���3�5��~d\MhD������tKs1<��_�@X�Uۆ��w�\l�eA)T�ݩ-d�U������5Ogx��:{�>�W5`�@TC��60�9���j�	�H�-۫C9��'�7����Vn4m!C��,�t{ܽ��X��:�O��W|{@��^�`��(���)�/���c����e���fW�R@��?MF�
"Xw���U��(�c`���<���Y�Y2�,��P�@�m�dB������G e����F�͘Zھؖ��qv���r�T(~��}F��n1��C2\erFM#��V>��H���d�D�;h�}2l5j�{��*>#�A	�B	���^��(��0���~�@+�1�����V,���B�g;�1[9�5ʵ���vI]�I~�/Rj^BV��/����/���EX8CX�R^U��:SPH?�5�'��R�b�ȵ2֒T�ϊ[�E"v!3(�ٯ���d���I*4XH??k�N��Y�U+�C������j��.�l~O	!��QM�0[���$���q�r���|�H�{��q���|���&��LV�D��ݯ �S<�O�X�T�mIq�Z�.7���d_:]CPp0F<9F����ݛ���	���T�#t";�|�id��B�BO�;) �j��)n/���ΟD��� ��%�z��R"]1[D�_dQ�K8DuPsh�(�m�u��4�� ~�Ϊ���)�{��T��?�G���=�!�ԛzYH����o����0m��;��������<օY	pʱ��׊�p����.oM����6���J�Ҝö�]M�d�̞G�J����p�@���oe����R�h� K�i��]�̔�z�j��>��2�� �Y�t�aPMM�%	�:��˒�,�x�\���-����o���4}?��? ,����9(!�{�W��~z��#,%="U&F�0�v��L�tN1L2f�h�5�#=���V�ۓ͊$ć��-]N��N��u�F@];�xu\�v.�V���Bu;^+0�6�v
�/P���N�.�=��n�?B�`$�c��<c���$x�]���.w�u�S�wI����]�P�S>���� Y�!{�]�Gvb��
Bu�-@���Q]��|P����ɑA?��GY���n��s�)B�.�*�s=�y#�����4���y�$,R��s�&�=W_�;bo���TR��GsH�H����wcT4/8ٰ���'fBs���]T�<m�XKj�C�
3]{�R���L��H��ӥO	�h�j��Z����1����S!���l̛��d����1u��Kv�4xI����\/��7e
P_�|�#�������5�}�mؾ�ja�)�=��B��V�HUC*�nEv��3,xN7o�ѥ�`�ѭ��U��<n��%��Y2�'���4����.W%{���Pc��>7��B���]�� �@�W1#۶K�J��^�0�����	�R���C���C/dW'� �D㶅Mp�zTuݔ]@�z��^J�|kX+*Jq���NwKc��'k�"��e��v�O�g����Ϥ�{��,S+�ӿ"��e�s9�m]$	\���M�����9���
%�����L0
sK�g�\�}��L�G�Գ"-���.�Tlc��8t���/�%��;1Hx%�;Jp��A�f��n�^d��,�+��E���+�c�O���;\������XN�k�Ȅ�T]�v-oF&�j뵴�Ϣ�1V<�p�S�88o8�k�Aҧޚ�Ó�^c��z�KL3��Y(�WKoɝ���@~)z�"u�����/�uYda��w1	�����m;��?V����2��'WҖ���>oln�`�_�{��S��
��*���p7@�l7^�3}�Ś7��j��m]���g��M3�Q�)3;pp+&	K8���Ҿ�r�,�&:�O�s�3���<U��F�rtu@�_4�䡸��	�!�����J�Sq}\��� ���%�Ku��M��uMk�W�A�
�&[��M ��ӰW���f���
cmT�V@�vU��Ţ����ԱiϾت�#�<4!�ȋ0C	�����z�L�%�ęC�vAAL�}���3B8����k��|���bx����p�c�#_��=�r���ٟP �59Rq}ok���GeJc7�I��b$�
؇O�N�k,�Yԏ��:}��U�v�LM�>|���`g^#	iƃ���^��c]-���ni2��[8yZ�t�o̽F�&L�n�߿�G��`݁r�����=>�,8�o|pl�ώ�Tp���W�����>��z�W�gQɋ�u����ډ�o�lm̑%�%a��|@ڀ��J��4�t�P��l���gNM�|�)�&��f"��J^����G��Eʻ��J��E�G+�ҥr��%x����0��Y�+�������U�Y��پ� ��.�Ѳ�Ֆ�#3o����$�-�X��BBt�j��ÁX}�S$�����h��h�2$H��P�)�ԣ�����O	��U^�C�����C��fp@�GN�ᖟ��A��|Gzw'����:X4��S��i��z:z�BD2�n��N��\���oPJQs�������<?���L�F����fy���)� �BRM����.���O��E�P�՚����Bs�	��	�g�U����ԤQ[�ؕ�RM�.Gt���[�B�^/m�{���2�U�I��	��-	6yq���@��[�X�5�Ly�yK��N�W\2r��"��E?]�hu̗{�R^Ӻf�=E��t�>Y D�l���r8�4c���6/�D�=�S���t5`G�?��e��h�n�O���E~׳k'$��h��ŝK 杵��Fˬ���p�~�`�δ�OB	��Ȋ�ܠ�]ȼ�'?z��эA����Q}��e��>l<�D�����1O&gX��	�p�A.�QC_{����ʰ]B�P-���+Q���/�)��h|'�v��Y���M��e`���g���o�ɮ;Ɔ�uu�"	��d����ew��y�@S��&lD����^&���v��N���I����KPy�v����P!W����>�;	�*:dl�S��y����^�w)��C�� �6/�+@y.�`b��o�3��}g��r���@�5~`!.��Wq]��օ�G����v���-��ӂ_�:SS��i��8�R����{�؊
��j�K8��}�V�2k�z~�,����cE}o'�``#2�k@h}�kY�5I4X<j�Q7�m�����^�g\$�%e6���K��`�^6V~vn�g^�B����[@��>�P�� ���{�!�5�e�X(G��V
l��Ju��V��RF�����,��0�x���[�^���#Z�j��Ф.�T����/d#�N>DT.��x6T@4��ۈ�S�Vh����ma������9��7�mnh��Rkim�@h�ܹU�V��>g�1.�JՀM�z�IB�]���726�r#�	����kQ��%u�	�d�>����W��׊;z@Y����G�RW��.a��&&����SU=I��#�3��
~죽��)�qА�8�l��	S��P���WE9��i�/��zq���=�7�SY�W��w'��"���N�Z���VyH8n�o�s�ˌ���H�ha����O)A���t�J݈��|*�
6�ߐ�e�Z箻����B��F�e�xYC�����:��-��[�jA��`�7iw�.���X�N6�9��k�撱�+���}1_��i��|����	����]�K,v`X�S}7rm2�k��j�yu��h]�:��|��N���(I���j�QuI�C�;L�G�Ύ�f�uv�eʞQUS���U�h�6��l��Z%�h�̑��@!Ǯ{��a߻�rM�nwVa��-p9L�b�4����#x��._M�^��I�d�m��4k��8X�����gp+��kq��Q��I�Av�7�A�9�R��2��͝ENi�F-�>�=�=#c�7��1�F���X7�`�ky�=����3�}m���w[����߷��[�HK�R��_��V��P�'�-�
�X�WY���&���ѲT� ��
�l�FZ'T&#}ǧ�}TH����7I���\���a�"��a����S��`i5��"�����ՐVs%�R�ޏ��@Q}�����˄s&ֱ���6 ��nBҥ�ĭf�yeB�EPME��"���r)``���:���C���xҢ��A�i�
�k��C'���Ue���leyF 4Xf��J9���˨�%�ɹ��E�~4A�=D^�.P��	 �k�௿2j�p�먊�=��]�$�T��~ /m��-��i�f�0�ẹ�h,�f�4�*ʜ3-�
������A����K�+����:5��X��
�^\��������`��E�}/����df��t�T`���	dlf����~�ѓ�����RE�V��,/ǟ)y�I��TDy/�L���K�ܯ}�f�qb�~z5D�_��M�I���3:�}ְU�:�z��r;GύY7��-@���MU������}��X�F�vX�� 
���?r�n��]t=��-��1a�M��J}ry19�Y��{\c�]ޤ��鄣��Ǩ�f+�"��!#���ܨ���1�T#j��]6�T�]���}S����C� h�u��Z��vX��GI�`��,B�#rW$�_��l]���4��-���,8�H: �M��?��S*o�C��hn��:y�F�}Ѷ���'ۚֲra5r��ߧ���p�eՔ�d�,$�/7qЗ�ah�|4�S}���r� �:#��ٰT|.W�/���s%WK˳Y�¾5��������s /��!=n0o|]	!@�� ��V�r?�~+�~Q���-���6�Jp}���2����	e�,��>��#� I��J6c�Q�q�[m<
�j������r&�zX8u����c]���2]�� �x�ڣp'Jn'T;��l���ZhvÅ��	�b��{�GWFn�x M����A:#��돝ɬ�m�1��:S��s�o�!`��ƀ�/�����7(���i%Hb�'-H��0f�{��.��m�4$�
�v����^�]ǑX��gSwV/j��!��3Q���,�A(�Ι|�R���I%��}-�PP/21kc�u���B)�p�쨉�u��~H��F�Z����}�]Ɗ7��VT>	 ];�5>�$�$��aR��B�����mwqŜv�t�;W�ɏz�!nס�Z�UuJ��b��@m.BGr�m�,��E��ښl�RX�%�9�d��^���`�l�^8�K#��{��'���9p0���hj��
'�q�?{���o	A���!��Ղ�]�M����9ܲ9>����̢<���{�[d4Xk� _������ ~�c��@Pfѳ���5`�,��SO8��t�z�,�KN)�mE_�3�ټ�p�۟wi>:(J�!�wQ7`����;����g��k�F�%�H��٧�`x��*Aϭ5�b�H�G	�x�~R�R٤J}�%!��/�?)���v����ŋ��o����I|����4��E�	(���.}� ��qr�kr��E �e�*�oM�lZ�(#	Z[��Li�������{M���k��F���I4$�fhCW3'[%\�P�
� P!��B&��ok����R�-�����]R���dx�_UΞ���&x���y��H�Z� V� �ZI��(p|��!(��	�!��fW�a�"̴�g�'�ae�A����i �mT�,���#(����c<��{�{�h�A��)�Oη�pr���a�
'd��I��J(cg_�\Pϣ�C�˃�q����Z�` %�Ijc	�}��7�\��gFn��sE�Kd�=�Y�,����!H�.�z���-�2X�T7���5���x%��� �S��~������{�-��<=v��ɑ8��d{�H��h�ϲ��%Q%|8�I8��O�� S�">B�Q�c��~L�����l�������R�N���Ӧ��F��	���c�3�+w� ��X/
�����md��\�S�H�ЦS|���Ls��x:��8x��T�J`�G�A�8��VLv���b�tU�4*ꑢ��	{��
�% |��%;�oL���=@F�����I@�����,j&�D�oK	�X�$ڋ��מ�cNU�U��|��/.�)�]�`� ������E�D�S�c��݊Y��n�1"�ߺ�A�����d#`X���j/�³Q\�E��=��$�(]��a͞���;���|��=໘[�`���g����ꜹi���r{9@��q�d�}�#vʎ_�J~�l����bv�]٣T�u��t�n
>�P�[E�h�#a6ڒ�Rݩ�\sn?HX�����@踴��B���Pr��g��e����%�sOp�z�CJ;$��勃
">������BI��vGk�[�n/z<S������Z�u��R���.�`;~ڮ�*�4i+w���)��B���tX�p�Qk�]�|����f;��y'���Q����3z������]�6�͓͍_���R��'}�k���HP��y�����;�i�S�x�==�V�!cDi�`�[�H�F� � ��ILW���L��U��:����蓗^ #Fs�U�n�+�5�'��^Vb���)���ŭ�k`,� ��kUC�N�R�.��D��w��i~�]R���U��V9�dp� w1Z%���K�޵�4N�n�g��$�kA�>%�xy�O������߃�2�9��n��P�ʎ@�I}�Nu$��$}w��py��A9��=͊�h�"�?����#�b�?s��ݏ��=2�M��L*�7�/�?�{k��Ƙ���d!C��@2e���"�jI��|�P���pu��cf��W�!�7"㗯ֱo����в����)���B�6N)���ٜ�܀�Z73�{�M���!�?����u���bȾ2c0_y�Q�0�Oc�:��7��\��&Ǡ�	F�����հ�"ˌ_���m@��E���
��3�����z@{��Q� L��RԔ��s��mC���{=�C��W�d˛����W̓��#�{J��"�o��Xf���JJ�FJۓ�WxH��Zv�tXD�Y���Fq���ԑ�b�<8䇘��_Y�@�XN����39�n,<���C�w
�b�N��vwO	�{7��)O!�1���$g��#}�̇%�A�Z���>:�a zCz�=d�ϱ��#;e	�Dy�fgM�b��i�b@��J v����r˲���hr�w��z�Y�,����KG#��3�kB��>�(*u�h���E�6��i�J5�	��|fR�>�8JD����]J�Fx3DO�7ŵ�%mm�^�rR��8f��Bn�l���ٝ���։��v����'�
,Z	�U5n4�!�`8��Ȋ��G�u��7Wt���LW�n����E������M�Q'픀��n*�v35���IMJ�i"�d2{p�����0M�:��l����ۂNL�����r���Wm����f��2;.]���TrA�й�Eh��wL����)��rnb�OTm�M�e��r��m��ʡ�)����F9��%�$c4����i�<�7�ӌ��sZ>��(ԩ�Yl9�?c�ʝ�)E��kz��[�*�b���m��������(Ըf��t6��h2�𼊹lb�!�2�)H��ĴW��t����U!c?��&ʛ�C�c�Z��&�kR����C�!@��?��]����Z��h�txm��qqܦme���?s��(�&v?���5�{-��5"e,0�1`��al��5Sa�c�ؼ�G���7���@����X�w+<�[�S����0�6g�^gӜև�i�l���<���c���V��=�P�ψ�6�����Lm�V���Hd�����~�5�����/{!�Lq�L)�6�@���A�n����p\��v�;#�b\�[����訶�V��me��T�b�_V�1�`���Pc3��d}�f|�#�,Qdˏ��XI�8�FG�Ն�i?��� ����=�������5���ڲ�O�*��&��D�qGY$����X�a�r��/�����m>��s�� �KSQR�I-�)
+�{4;��IՅy)� c�Rڨ�K\��n\��O����r'�(�.��ul�����@	N�<���$��?���M`{���Q��9�y�)�&��}��X"�eӂ���:R�u�P���h�]:!ЈQyu�ĭ�<����Rf��i��0{ٜD8�_m�č��g�:#.�{�c��ӻ�:#�A� �#h��j��l4�%��솕���:k�g�H.Գ��ü��c�,ɫ�)��2�u�3l�vA���m[#�[��gc�}J���g�F�(�U��4!૱��˲rJh�\h���S����L�Qk`N���YǢ2.s������۱�>�K���0	����V���+�=�{i��4[W�ԛ���M� 3�iN��93�o���P������b��b��҇c(�?6��*�Z�M�
Ɔ4�P}�jD(��CP��G͊7��z��m�X�OӼ�'�]绋r ^����&mh�%��R�1$�9�P���i� ���x�����d����@��%*9+T2N�υ�Fey
��,�+:�o��l5����C]H����]+�ᥤi��1�Px���maf@�0E��rP�`F�`=��snًZ��l2�Iڃ��� _�]�T�.�9"	myj�o2f�s���T`$Æ=�)=��i�&$涊���{L3Y�������%4x�t�N�_���1��t�k}�E�0�3Hx~ �{�;�}�'Ю�����wt�q���|�2:u�l����|����0��l�T��\h�����J�|�v^��^AO"̕���ܚv#�=���:���ǌD���aei֡���2~(��ҬJ$�'5�̼��e�%��H���s��|��#��t�N�g5[�`!]A�Kw�| :�����	27B:m�$�S��z����u��_yq2����;:19:S�f��ʘ:�%#k-��~{�ېN&�a����v���Ԛ���k����kb�N��72����Kѱt�^A��ޜ?0��&��� �H���Kv����� ��^2{�Qw����^�;(��bK�
�X&.G������\�wYs&�&[�0�W�>|Xz�$�Xz�е�t���n{��g0��x ��R)�T)ZD�78�:A?��p���:f��{��T�lSWmu᥾�-�X�e�}H=t�f���`����{C�0�GK:��Rv��A�S���0�+ڧ�j�R�ea����N:�hm`lTo���k�~�+�dh�QJ�΍ ��<�"Zb�� �6{>�y	��Jܬ���[Zt/a3wјu��� K�b�/Y����e���j��8e����g�yѩ��DV N�G���x���/�������q�:�%r��{ $��P^ _I�3�c��|��Q���Z����uϸT���)G�"xB;��������M�B̂������5FG�v�[	�y0ɒo���uYj�KE����0�U�M~��&D�}���)��f���Q�s,�ԙlf��l7A����:c6׵ޞmˆ�qT�r�:N�0
��۳�=�">��U��I+�5�垇>��ږ�b���Wu��\��'v�6UPs��o3�rg�6y_1:*-��=�����r*C0��x��s��S�Z�PP��J�[*Yj�B���پ=(f0�$�觭��<WL��cT�:ۉTa(�VmdȔ�,��/H�˵(�cTm�y��Е����0	郆NI�v�i���s�x��!�/�t&��a<�	-���x���e
&w���]o�,7~,C�V�w�=.-rXP�F��S��V����˺UY��N�xǺ^E��L�#%��e����L�ˌL���EXnLb:/:Y�媷�b!D^*q��f+��������g�ӹ��z�ecz�+�»��`�-���p�\���Md�Wz�1~O��$�1�e\���p�ɤw����!�=h�ڄ����'w��.�e�b����ի���mP�!1j�y���7|6,���/!2���;����~��Y��a���Ouu��U�><�k�f�b��ag���P�0�b���B�If��ki��6����Xŝ��ىbS��8t�E�ͯg�<[���F���)� ��ߍ��}���q��Vd7�Ł���:�$��a`������8�q]G�r��Y�p	G��uf[#��P��"wWGvd��ZRv.�3'e����z��k̰��ާzY���9���j[�MT`���9���g��E:��sB���$S��,\����v"���\���z7B�)0%���� �B�@��d
J=���o 눿�4.A�Hk��&A�t���&�4"G7�(�b1M�^��nL�"�x�Fo(������=�+<��0�:|�ɶ��r�m��/d�Ϥ8�o�*bQ�8�FA���_+�`\����<�C�=��B����CF���Ͷ<_=)K��P�m� ��w�<�#o�~'�bI����;C�_��`1���*$#��'��Y��_3�����]�Mq�  �9=(3$��`3��>�Ql�	�?m�A�!)��^����4R�9њ�k.u��K:L��c/���5T�Q�o��T�{��_�ҬA�h
��_��8�
EA=��%N��J�Rs��q�C��'��e�S_F�ބK�#_	�{��G2�D��uJ���+Dr'	�_C B6�7�mz:��^rɋ���b���3/�8ǼϽ���p��� ���o(�-1����c��L�a�1�����]S5S��?T����]+o���Je[AYv;S��Kם�6_�����1I_cr���
j��+*8���<��Y=l��!�?� 4�#]�,�U))^.����x	�{��<����ݸLV0!�P���R�?(��@k<�d��t�a��_��|AE�E��0�H|�ppa7�H5���u��!�XT4ƌ��&�_8�Kƥ�G�?�_H� �!څ�C��>����j�⁕0�X`���#�8���<%v�k����v����RJ��g�e�a��՗�M�O�KE�f+���ph����&o.��AO�8���\h^����^Jf-����-���Xs��D��i�.�F����͍	��t,�.|���N>,�����;ܵJ�z��6-2�J 7N���F�m�08�`�MW��pW�ϳ#]i9����s�c��{���#��b=�]�U�鵐V�^|[d%�%ak���&�ay}s$(^k��iOaF�h�J��fS���2�`N/�k��+.�C�t[������1ӭuWa��G��$�x�5������8
�nS���A8��m��<q,�������;��l����ƻo%�aaa\��n{�w�K[��N:F���/�y���ou�da�M�fv�f��`�X ��V)*^
T.ǈ��A-'ɣ&Q&��8�̧�Q�>�=7pdШΚQ��=�i�W��A�r���������)<n�AUm|�f��E�{Y������ �PX!�f*����y�B�Q��a��2$���i2bQ����S+Da6�s2��h�e@��cFs��Y-�o�(n�aG�u�=������-�~�X��2�V���2���=��yu��cm#�5��&���?3Id�2�E>m�[�a�߹^�"W��$٩Wv��E��K����(�`��CNsu,a0a5ϲ�^����s]�[2��$� �R¨�hz��J��j�����vDS�F�e��m��㺊���``.�����*�d���-���E3Ax-�8lwC�$DJ��T��,�=�'�$�a��^�3�����ڮ7�I�_ �c�u�X��$n/qW�YF"�I���y�{�Ҏ���8��а7������Hl�$&0�)KK�}$I��Ïm��3�Hw�ix�*(v9�����c�ʺ'�I��?${!yd��R�Q/n
�|ڄa�"�?gqO����4��!��NW�2/�PT�R�ɬz<J5��Swc����e��A��^��	��� ���z�,�La����R$,�� h��A�/8N����-S��O�p.J� [Z6v��eAu$6�U��q��_�zq��K�-G�Tk|���;�^�c�a�N�Dڍ�V<��U�F`��nBE<��:s��P��f�8�Y(�K8iH��ӱ�E��%�l���	q�ϳ�:^�4�3���<��%V���Ī��93�b�Rg
4�9�j��������l6ǞZH���/�^���!#l�Je�������l$"�G
��06�ւ� I�@�øBwN�_$ֵ���k ���+\<A�Tm���/s|��T�b�M�u�盭b�0���淉QP�AJZ�/Oq��}��&���-��׎Y���5@��6Ǒ��;5Ǆ
�7��۾��EӰ��3
��sY�-�@X«Řq�^K/��bv���cm���+�lp�j�+��c�>�V � ͯ�e����f�X�t��[��K;2��a���Fg��������"kt������K�3Q��qp�Pz<J��"��v���T���I�e����7�r^Jt1+@�r0�v�ś/��m��B,l��ݶB�����P$�xX���� z���At�+����h�V�`zKJ���C�7��Z�.z}l���D����[F�CT;�E�Y4�����I�J�� �)��t*����(?�HC���P4���v�*R��b�O��0�r�mk[��*��ӎX�-�ݨ�]�Q�y&z�4���?��urݠ�8��&;"�u�9����赊��u���T��IMs��0`�E�1�62Ťh%pNz��>=^R���$0�n^'�nH?L��
�^�R<��\�( �� �4V�_�B`�l��U(���ǅ�֪`z�w��E��R9��qC�e�!~�.
��ζE��)���sJ�s'I�Am �S\`�"�ȯ '$N���AV������!)!F�> �T&�I��0@b<��O��)��"R���Z�/����C2���E�^�
�/�?'��@��mݳJ���̼f~wϰ\\�����t	�y�"u�<s�����	��
b��v�M���s~�!=f�G���+���=��S�²��!u�6���)/�%a���M?������bB@{C=pIf	�U���Ͽ��4:ᰇQ-պ����=��S�cO�p�昀EhtD��k��TP�P$�yQuh��K7���)�7���3�[͑��k�?�J�Р~�B���_��t8�E
Q�l����[m��"�EJbh�r����߆/���> p.�H{.[.�:ӯ�����V���dN�A��f�ٱ2���N>�����ˠ�x���v�ڤ>�pB�-�w)������k�1��Gw̘��_���Ͽ�aU�>wWk�=����ִF���RE���Cj�ȫI��Z�l-0�@q��{��5��$*[�s�j���$�l�y8��@���@��>�(���e?,"7T6e�����:���&���G���$MW3��.\lD��C���Vt= t�0��z��7����6L��LҲ�jǷ_��@N\P�;�;'���8�b��[e��H���e��ŭ�5r G�*?�ˉ8aL�n�
�t�j�����*o_Э`د?	�0��K�[��c�\�	�.s���h3ü��$����ۻ/�7~T���4>sR�����c�޵����w�l
�Y�S͜{�M� ��{�����=�j�~�R�w�ii�f�~���q�yJAE\�_��M8ּ�!�ImW7�G���ZJ�N����3>D0���Z�x� m��VV��_�1�|��$s��������wn����k�j5�ʀ�2���â�	�l�q7)�;�����لڔ�*��N�. 65�z�?�#��n��
b�/T�)(�KL�����I��n�����,�Q��y��om45iKV�2A��M�bK���c�＃8�,�(-�s0���UtR-$�Xٔ�ۜ��z�T <�o�&+r�G����_��/H���$�gx�i��cK��b�/������s��,J�sn�x�H9�Ţ\����$� �1]x;���,��[WS�=2��%ݟs�5%n:Өji9����Cc�
��u������E#o�d]�	ԑOw���츋�D�GsH�oz/z��2 �F��on��3�ԖM���J3:1)�pxO��; \��O�_fǵ��YǰMp�0�k���%C+�<���2��\5�[����P�O�]��uM�dM�8�o"�^r��2�ͅL��g��h�d��f�:�t��z7|ʊ��6�kl���k�6l�L���=V�|�|��8�ʕW���lՒ�^��2qO�n���	�K�����`�|�\8gi8� ���M��B����␹3V��H2�M��Y�ÀA سXvV��c�2M_���eӝ��ڪ��b��u�0��i�w	h��1s/����Sv�n���;jW����?�}��4k���᩺��#���ԫ��Tv��}$�x��h�ˤ�k��bj��������]��7rn�Ɗ	��o��!
�m�I���P���IF=6��6���B����� 9��S���/~\��&l����?t�*�F�Gx=�$�?� ��HL̚��������44�1�����Ɵ��l�
��-,9!�	1��G�Î�9k��e��G�ɅW|�W���]�mw�0� �/�0�?�����zJ�˄L������6%�&kC����#�9"T��Go��ba�`�gn�Xm��x�E�à�N�͒~��(���a�CN�����Y�~(�%jh��NoQU~N���M[��}��p��
&��""��o�;�ISgv��l�8��&���� Ώ���<�,��< �i��sf��O���Ϫo<n��h~�Z}oqM<�y�Aƈԣ�w���W�a������ZL�����Ň��:��"%�Z��˥Xh���Kpy�,Nq;���T��(I ;O�&�^H�ɷ]�G���E�̅��^�����x�q�OP�Ӊ�`�����=~#j�>�������� ����y���z��)%��q��Eq�&��`���Np7�E��j<i�94��Q��G��-@�v�M�k��4);Q�s��.� _q�l9ԏ��$0G��J�v�e=�/�@)k5b�q�#�H^6(ۺQ���bB��Vꉐ�F�&��d�lЗg,�Fh��	��A88���?iB�Ћ*�!����	`��ܒG��:�2{Rt9_DT�BOȻ-��ٚ-	�ZW4A%���DY��������S�dl�����R��!ʛ:�ȸ�5�q�j=��z�(_ D�
�\F�-�Q�Ua y�. �Kun����:˝Uč0i��9o�1�O��\�&4�uxLX�ٿ=H�5���ЃSUn���V%9��2� N�:�'L��C�/�dJ��-�e�T�,ӷ��+x���r�����*.{dT�����D�9�����(�y��J�*�a���d�\��F�T�mi$�=Ȋm鳬`o]��]��JiS��($��D�ح�*yh)l[a2��E��O�Q�)��v#�&���̷`H�X$ ���������3�8���ݲ9"%�����eQ��&���z�h�O��<0Z�+�	@}��ڵPaQ�o�s'�x��匂ӇQ68p.�*z)0�F�K9V�mO�q�md�Q��R��ȣ[�i���o.���P����ZoU����lNqjT�����:>K�4�:�rι��W#�C��1��P/�����f��q�P�X�43��O3 E��0�k�s�����G�i��μ��s{�����tV�ߓ��4�7�z��'أ��	]�`�(a�|�X�]��M1�h����ԏ�y�Im_�zŬ������?7,�έˁ�5sU�Z����8d:WŁ�n����2��.���6:�]�\�I��4�}ݻ��j��`S8p����[
:��'>�����A}�
����Xfl��Ea�gi�~�ϙcӬ���[�益���e!��I�++ƗZ:��[KC��|��Of�0&̽ï@�ߗ<�k�h�V"�`��@��M��i<t:AI��CO<W�ء��My1� *H[�}��|�����bm���K�Ǻ�3�)��������Z^NY�}=KI����ٛ���3#�	nq��yj�CHn��ʽ�S ����u���U�Tb�TZ?�i�C�&�3M�Ř������2>O�XѫЃ:-��m��{�.QE�����������9��f�G��O�]�[���y���N��������j��b.�����L&�~W��
]��hoܳa���rS3Tq������3j�k�زi|i�FL���q���L��������%I{�<`����*Tqd��۬<�3ݬ,�l����p$O{<6�Q�Jl`.U�3`����!��7f�+DZ����D�k��7SЮ%8ʖ#�n���o)�Y�Z�i�Z��K�IF����ŀS5�����`$�n�4�,ϧ��V�;9�kdI��l9�X���V�'M�Q�/�����[L�PLk�>j�zG·��ށ,G�n���{UIߡ���-7�j(!��H~�ȭ=�5��Y�'}����K�0� �l!�=��Q����p�s%,j�Ř�''}Y���Oc��%��<�`��A(���
19��Cv*a�՛�I��8�c]߃r-	�����ƭ����`4��*�������@� J���tv~�2�����˺A=Ԕ�.���V��-u9�䨛��Ԣ����`��!���6����7o�/%����8�S	hNa�O���
XB��$t�d�<�K2`�K�����P�_dPf>ԕ>���mRB����,ȶ�;�Pjg%��.h�|��Ĳm�]���>)a����ý���5��
�w�Ǻ�.qX�!]��ݨ,� �F�]�@�YXW+q��f�_���v���|uV�zz�2��ˉ���Ix�4ׁ�@��v5�gd��\(���X/��:�K@�����w ���
\l �9eEc�V�EF�f�)c�j0y��!�2�����Ëj��Y�B��eGD|��b��V��>����+b^\�M�Ɂ����ZΙ��*�	��6��q��8�2�_�̌�y0������_���U>��("��M#�
\�50��ng
�����7�rI��*➨#�k�D=��&�j^��(:�:���/Y��l\�͖CJ8���ʾ��l��J�E�z
BI<=���I��\\h��͐���Y�'[�䷑/X��@��g��ʪ)�z���-s(kz8�<�9�sI�@2��#P ٨.�+�.o��kS!*��}�%c�&#�������Ӓ�2؄�9�l���C�m�'����1�"9����-BS�F��<0�#�>1v	���[	�@ϡx�ګ�r�FEt ��g�p���	uco�,W���:N�qO�Q𗞄�_n�d��³}#���	'�k� T��:m|���}��\�~��e��SK�YqDH^B.�I���R�$p�wS��
�}|�=Mje�zY�9�y �Ҝbp�4+%)��^�Sb�q;�u���9���f�����@o���=���������t� ��Ա�X�Ѩ� ~+B��tٌ���'C���l�4�.��o7g����b$���������Q-�F\aSw����g���K�n�xU�4�؀�\2�+��_s���&�D�"`%�ݵ��j�[.1��n>�ğ1+�R�P��A�$xI��;�{�������D�U)�'�Ē�D�kc|;+&���վh�*jI}<26�{�Onaf���P�<���ᱵ�3_�pnDT�ܾ{S��L��7�oH,��6��`����hZ�>X9������t�d�2�K��#�����f�4�}�C���wwB�Z�e�W93��A�=ڤ���XV����8�,$���#���wTV�tۀ趵��#8Ѐ��b������a'\��!W���ȳ�^�<��eG���/VӋ�U-�j��F�(�1�����|҇��Oѕ�:�i�)Ɣ	��DΛ�W�f1Q��g�&��Ͱe,[�����C���e���"�{��;j�Lkd�.I�Q�FDdX-Έ��#���6{�<0��]��R��j���5ng�.(n�&�n�0ĺx��J��X����? 'uw3��^��R��lFu���Z�:���P�b���~k(�rz� W�Y�[��RW�r�c#�?��ӗ� 'n�|�.�V	���O�n�՜���(���W��ٜ�#.'�d��7��H�UV."i�� �AB��ږ~�/��I�vw�7��su^2� 0g�*��,'��H1<��r�%�R[���$�~Rg���^K���o����h��H^=c�d��P����~�����Y�:�w��O!:��-Z�����Ԭ����T._я�?�z�QtI�^Ԯ�7�8O��!�)[��k�.;�`Ҥ����#aͨ��|�5WnPO m��=��)���q�UƔm����5���u�\�C��U�u_ƕ�G��,0j�}�W]���Й���'iX|�2IS:R���!�ȵ/ԽR�{,����G�]��m:����a1J�|:��')&�!�YíB������c3��=-䳺nt���H%DH2b�u�?��ڮ(���4G��K�}�{a�OQ���G#�u'R�8<=3@�E ݦ�Ki#X�2ᖋ�	��1�}7����w���m,�-��2���}ßb��*Ev���U|�Norf=9���5�S �u+۫�˟�x؎l��L�-�G�B�S��w��K��<1�io���Ӄ,�w��,d����B�|2�X&'�(Q?�x޼�~� �{H�.f����;�f�'z�v�b��&�"��9��^l�4F,x=	��� Ǟ��O��V^h����ڶ�u�l�����;��n*�b������#�Z/���"q����
�^����S���Ȅ�|��A�j�ױ���4�r���J��^�g�V}>��tu�o�5B�_�R��c�BW�^Y:!`��_��_/����S~(� �|`�˪�Z�/��y,F��Y��7�K0Y���"�b�d��'��!M�ކ�����*�-��zRɔg�ˢ8_��Rk�5Z�Ձ����������\��Wd/_�d�˖�"���-D1m�<�d�q��{aKmd ���԰p�=�n�}����ii:��ǡYtql�/=p����]��]3~�F�nwj���R�����=�d�`ܙ2K"=�p���~�������v��[>�lo,%~��%��{��M�@�_@�{.����F�V�����[^�&���ϳBv_<ڔ��(e��H�L�)O�&��;�r�n�Ĝ�|�>�c�
2��Qڼ�n�[�n�ܒgp���|Fek��C'��s/[ ��ZAч唽Yy����<��ܘ{ݜS�h��2��k�9N�H:B�ˢ.Q����g�ab�I���굞���>P�H����3[�՝Ͻ�e��Ej�߄=��ٮc�n�0Z"cX�Ԇ���_d2��K��M���:P��z�9�� �LRj��:-C[꺬vy	AoY�8"��	&�\�cV~�A�è�υ�d��R1C�mk��X�䥳U���qG�"�*p̴�r9
�]�a�Bޅg��>�qP)v�K����P�����%�)��=2�11�=l�8�M�:�V��RB�7V+X(jk��1(Z�LG�"�}	��-����1�s�bJRQ��j�;��R�0���lږ\JTuç�ܢ�RK�km�㗡_�J�y�f�x���r��֫J�݀�kTLQ������#�3$���Y3�W��&�^z�����#�3ϣ�_�A~�b�Sg��uGI[��@����׶E�&GR8P�{BuEۗg�o�ʮ��\��yJ*����;���:�����#��l`�(�߽��?
�}2zH��==�p�Ў�Ǹ3Ȃ=~y$DY1��)�W�Q�x�6W������%�Y�<����lG�L�O\Δ ����Ӭ^ɦ���2��[�M�p��J����͗�UF�gR�BZ���?:���3��v�X�O(?��c�a/oy��W=M4x���C��;�"���ǩBI9��\�a���V�=+�J�aZD/3�D�b$G0�����8���%Ŋ$�ڨ9q1��A]'���7�7Y�&Q]���Zo-h���;(���<4���2�>#�"�
1�s�y��M���L��}�+\� ;���0-�c����g�@?�{�E��0iQ}EZ&T#C��0��t�����m&܅�����|�?�?�(8�9��Z�ڸ��k
}��L1�p�ib�����e�P���qPS#��2��q �"�g5FoO��|"�����RO#�W���H�>��0����v��uh2��x
�@l�"uc��fcX^:��B�jo���Ej��bGձ���7���Zq�ZՁ��@��]����U�� )���3h������Tt|�ϷjY�5{]�W5��O}~ԞJ,#�o�͖36E��[��D|Q��͑;�߭��ߘHV\�6٭��I�!C��(���x�,_H�FZIX�>6�e����7�P�$uE���
xu���M��G "��s���<	�*�%��fT�@''����I���Nt����R��e|�G��V���WA�.��ƨwo2Jx�aֱ�N�i,�.l��2��td���L�դ;���u��m���}���l�o��1�.qV�w�w�} }O��_�L{�q�s4y�L<��!�:1tؤ�d�ab��d���$"4S;N�/8)%+ߐ��sRM�G��dƑce�+����K�<�@�8��B����?<���'�Qv�%�zO=��B�
��%��(���^Z:~𷳛�ӛA��ֿ�� ]��Q�G�>�NzΎ��l�w�`,ѩql]6���J�G�V�O��`@���-y�d�G�-I�%K��
rz�,"���}k\M�W[��ֽF����n8>�Htnq��(T�|��11��E9a	�����b9��=dЫ/�܀�j�~�1�ɻ�u�,�?�?�������|G�Ԏ�݂���S����}�2D�Ê -���),,�`�+i��W<���G�lyg���jmv�NA�&f������>>eќP���w٥��5��Ԫ�T=K��uS״�N�W�$D���$��	�΄o4��`�F%��%}�J ���sW�@9&3�pԤ/�-��LdڤQ�_Ir�D5%��6ߧ���8��D���;A&�[`�n=*�-g#��ZJ:&⢺,��S�27r���J���`�((s�iܯ���(7t���*4&z���r�*����Ϯn���a� :ꌪ�(�Q���Ren�D8)��Z����?|}~�g�.��������ّh��V2�4Z(�=�r6Fn��Q;�p�`YT���+vܖ�<�x��3kaM0�a�מ=wڽm��͸��C����6i�����fI2�u�q���2��Nw6�z�0w�����Y)�.���ʿ�S�7��D�ld�M>�/7{�^��d��6S���>��SÆ�q�g�N���?X32T��+5v��g��51�Tn��+L�~f��|
��۴�d��ع�;�ZS�@4�u�!��v"����V�qS��x&6zD���L��{���͵�5�s�����4b��=͒��Z������?���ʛ�Ma�AⱹjEqا��Vh �vo�3�&C�}V�K���n��U��;"�Y��.�P>���[�qEVaOΘ!�T=c:����E�?�'<��p���0�*�iJe1�`06I��s ^{��e�;ù>�b̤8��p�	#+���2~L�%.
vR�E(��uK"Af��agU�&���Q�Qqo�ZTyWYn�%�J6FH�}1o�-^�-�<W2�z��:u�ƥ��[Mo��¢e�e��#2�kkj��[����	�Q�>}:`x���!�?PO���B��k���F
�� ���1���li�$���A�����*A����b$Я7�����p�Ύ���L����V$|S�q3�wr%1�Wt�Wg҃����D�&�feT~����4HS�%HYA�qU6��@$1X�EPm���(��u����e���c^6���ԏ�N��H�~-e�մn����(�E����F ���	���E�?W�uq���
\���Y��Gf;	i��<:'#oޮ�<2�K@6"���ެ����b��(�H���+*��h�eZ�it�3���ɻOE���Ո�{�8O{ɊU�du�5a}g?�zO&qw1N�ȷZص����G����BP
8U '���]��'�Kc@��	�����v�Z�7dw&/�0�2�fР�e��۸I����6.�A�9[�<Z �v�M^���}r��,9`W��\Ӏ���_'��a�"}�y\ؐ���g��Kjss�YU#��S�c�F��qKDq�i��D`H������V+��9��8ڂ1z"��w��YT��ȠH�i��{M�Kf�E�%���X���"�'V�:���.����+1��t[����__Ҷl�X0ᖵ%S*P��r��H]&�^/��M���r��l���-\J��n-��pS,Jvy��K�a�,@���{���oY����Z�
v�Kk��o�6���5<ll2��X�^o"�
2R�4(|vZ.���.�2'���s��	m�R�`�˺ �g�-j�`I[e{�ĐC���3��$E�|֥�n���bȫ�j]=>���U�2�lHd����sa4^���ٹ��rp&���������y��eW�U	��3Aܬ�
�?=��y�.	��>�nb����Xw�����I��.��Io �3�ZBq�����M�Y5l�:b��BX��g�^e�鐋:�Vĳ�t �w
@�1��C�uIv����%�"���]�:��;�#�{�ޤC����OL76��'�^�Qi���("��b��A���Q���QֶD�Ь���X�u�z8*=�ǅ�a՜�N��yVl�Dm�G6Nv �q��` .`t»�	]�3u�Ӈ��͇�!��Ż|k}vď�ΰ���p�;�QM���i�
�WS�l�~jyQz��h��
�g�	�*�%�H���]iΪv�y_Bw�=A1i����y5?ٍ����3C6�'�'t��`}b��gV�2)b. �C��,1e��-��+��զr���Ru�h�!p�9#!ҿ�
BfU�c�:���u�c%/ �5nĠ��]}XuTm?r�e�̅� <��1�M�����ߘ��-����r0�oGt�Q��|�4A��=��Q�&~
��$���|��T'K��E�Wh���F����܄�- �x�z(͟����M�ȁ�=�/w��v��Xz��܈�`���<xo����|�Ø4A��b�v��H��5Q���%7�Q "���r=�bsy�<���LI
��"%P��pHH����CN)Ӊ���il�V�ZG/b��5�̏�i�=K<��9���}���[+<���&ۘn࡬@X4,PAt(�=�i�#��Y���6�#������a�g)�`] �ѷ� DXS	XZ��r���6���Ecp�̱��LQ8����GB��9����O��As�1Eg� �~8����8��+���nF�o��iם4�F�=�].(�ֲc��ɭ���+�;��Cs��+z:f�F�D-�y��%�[�+��z��y�= Z�"n��9���9u�>h��E����m�q" hR\Ȝx���b<?Si5.�µ�Hތ2��TCWI�Nj��7�{�ҏl�4��� W��,�Yn��/�4�)9a�����\[�6l�S{�:[$#���Gm�yX��0@���`9,2����Y߻�l�o>B�A@�ܢ&N;���>� F�5;<��tg���ݨ`HZX�p���j���� �mRU2�dJǭ�镍(I�g���I�>�:�߷xq#��!��_�w��%��ksL�3���N�kR_����s��}I��b��E"���DR���S�E���� ���k�l�Ѹ��&�c��i|(���P�Wv���d@����lq2�~�q��3�[j[x�{W��7�ی�$�ח]�pa�:O�.OҜ��� @'�skY<��d�3G��eS~�$Z]S���s�K�<Hӭ��iT�c��D�|�Қ���������]Y���q��<z��|���� ��o�&_<� �;�ye�T0|]�=���s�~��ZC��-6�F���a&�h��=�ꅗg�X�g�/�ϋKc��}����(��J�6vI�y�Iiq*����I#�����ҡL�P�Ǎ��4HF���Sӗk���f"�-L��J1j,���	���4>k��z�����J%'�TFe�xAQk�z)�Ll����	����}"�����@���TFSW�h27��ŝg�x<8�+��l��������"á�u��Vƾ��(nyh@��U{�p�z�}�yæ�CY�3��W�Y���2_�ѱo.���ƪW&�|yqJjWw�#?t!�^�O \"����i��*���,�t���CeY~*�?�7�;��L�l,�&�Y�PaT �ރ�K�z�w�9qH�h��F�[�I �[�� �e���0e�������~xi(�fw�AWׂ�G	��Y����-M�e/f�uT���E�:u��aNaBM|�֬�K8(k��<�~��z� �u�e�1Ww���xo�w7D��q�CL|�p�8k�;Tys���(�_Å�Χ��1�����h�$X%v�L0:�(�֋铐� E=]ė�3M�O�̋�\�q�po�*�� �>�u���ʔ�������1ˏ%�UC��n�D�#g�gF�`qiH�T�C��k��7VoU�)�r���B)u'>^����v���Ģ{��	b���a�_�7Hx���O����#����8D�ʲ!s�F`�HO�t�I�_:`Zg�cW_<�}��f]��2
@j�EP}}Js\?��Pz������hm�]�����15޲��+յU��Ҿ����=�b��ܮܼ,wCԏB�2~K�K8�c�500�s�>����hJ:[�g������>��CZ}!��!F2�a.N{���qS7�~~�1t�y@�ǳvJx��F,U`ÚV	PTx�i�q��g��I6l�;��v����$�&\��a��$l9\��;f�/�lEg����W��V�Ӭ��5�9f9 .P]�����W_%'�\a�9���O�i���f����s�"��I��\���Mf���i�X����B�z��9kA�����t]m���ͥ�	h�v�sL �Y�@(��q�=��?�D�9�$�
�RI@�*�J�1��~���2>\9.���`�0��v���ʣ���Sbq!K�ue[E^���\]%  c���N�:S+���yR�gM@9�p��ѿ*�7L�����C�Gǚ@h>8̇�JJ����G��[Z˨�9!Ch��_�y�/�߆;	΍G�X�a�ox70�Yu��m�}�hLHd���V9�ef��¾tnh��J@�ٴ�u4�!�m����x'�l}�Û|��!"�n���m�Q���w0���7"l��؅� U���$F�� ������������n1���ca�|�H���T���?3;,�ྑ|^
ں{��,Ļ���K�\��0�8s�QLd!b\�m��9i[��)X�j���ؠ�ƞ}���P�	�0n�AҒ��TdWm��-%>�^@�?
��P�n��K�%)���ܗ��DF�R�Z��l�G��6L�<N����$BC�Έr{0}'''%z�Qҿ�M���/xxef�2A��D���?�TO� �ǷC%���r��cEo�����w��J��K�ᝥ��zLG�Dٳe8`Y#e�����5�i޷2����1�!U�����ׁ�,QϿvI�c�_��6!)9؀�qjIqL��3~!� ��^=���&��0a�)�7��(C��-�:�*�ǟʱ����Ȉ#I���
ð)�k��� ���0���(�����N���CZ�EKW+N�X�a)w�T��`̎��Pt�k�Q���.(������ɔ���!Bm���w��Jˍ3����%�h�a���k�^�q�Z�$(2�������b�I���� ג`�a��Vaǳ\��覚���
��Sy ��vu4ܣ���I7��)=��p��:�D��)��8��y����L�J~��J�b{��N�׸IʻmO{�\ǈ]=���8�ޡȖ0��"5�ϸA3��Q�Sv�x��k�ʨ�!�]<}������ �y.M����T���Ә�Pw�c�NP:�-�R�GG\���t@`����)�|�}��Ϛ�������ު��m�����U��R��{�qM�O�t��> P�4�#�a��x�[����	�.)x/���qٻ� 8;�h�V�J����
Ų���]a�� ���i\Z����R��'�����S1�aH  �����D�v�p|�!�X������x4�Z��W��.l�L�B�!����8�0�o��ׇ�nt�䔻ǖku]4MD:�JƇm�2q��΂��dKz�G������`b=�X��)��#!~0%"�KD�xfK�;.�rM!}��K4�6�F1'�6���X��b�_��ϱ/D�����f1��)/p�9N~��I�i5��7s]9�k�	�M�}�l"nⅹ��J���O�Ί|LV(��+C6|dV -ɪ=��n���F�O	];���d�sZ���9��K.I�L(TaAD&����i����h<�X��E��#�W��	]��p��ߛ�&��f�f��O���
��8�)�3��;���&���.�n�=mo^|��n�L�a]��'�Y:g�ө�籷���B�xF��)Ks{���ڠFZx8�:1..)��|\�H��;��g���7�VM/s[K�8������������i�)�����VyX��[���$m���4'�+?u�'�� ������օ�@$���C�K[�qF*G�����hEkͤ��}r#�P�[%���w���8ҩ��?���K��rSL5�t��AB�pno��;o�\ѓbW���`�E�G[|�> 7Qu�˺'Ab�I�a0)�w�L �N�װ�,��X��w(��r��Qq{��_��OlG��y�޶��?�j�2�����u0�8m^��ԓ�Ȑ�ש�kE��g,jK @h��S�l+cTCMМ���%C:h�-6�z����DƂPL��g5�ț�|��������,N����{��2�Q���ժ8��t;v���	����~���sh*4nD��Ir�%G�m[��[I�+���` !�(�M�,m'[��Զ�bb7N��a:�Hi�^��,���?�y&,���� ���Kuɳ��b64^�>�&iۛ�Q�A�^�"�m���gg$	"�XGU�o(�0(���v�{p���~��{����������4Ё;u.Kkw@��(���D��+OwM�M���K�����n^'�������Au0���	H�s0�4[#��Ž�AS�}�IB�ݥ�$��q���MuF�ϻ(� ��5��Ә�޾���|��Sk7�w��J>��8����*��ڿAl����D��#�b���3�OuOu��Sy
�f7�jr�&�[!� ��E�)K2�{��H���t�e��Ԁ��@�}PMe�B?��(��}��e��P�p���Е��tk�4��%E��]E1*����[��4�_�~��-}P�'a�T�f�*Y�/���K��Po���?K?�����0���0#�+�1Г���C�Z�8��/_�.��{�ʯ��'�{+|L�	����Mg>h��v��,��ǎ޺8e��K�d�ʕ3�*`eb�&�М�})�M	u9݄BLd�[�p�h;��ݐ}�S�D��r��*U���!��9��Du*<�S�\sz2�I\�y.�,`1�y��jK4�R[�����;�=�L�$7q\c�� ��,l�F�\�)k�3߄��Uܥ�.�
j��6��gN+mlR ��ۂ���G��:�ob��s8�Կ�Zj��`���n7��(g t�z���5&�m.R>�B��t48�!.��C�j�*���̥ ��~4ÿ́�ߜ�h1�uQI�D�u�<F��D�tivQ�ѿ��q��Wh����v0�.�9�ޫԍ�M�p�3-b��"��$su��42�B�@	Ws[|⯹�i��5ӎ-k
q�0݃��zߌ��Z��h����H����t[�iJl��`7q�0J=�ZVT]��r����W�ӑ��H�08��D8�%����������U�$�?a��w�YǨ�gaӀ.?���Kz��/G��*�<1�p�˙���-�j:�N�s�}�Iɱ�Dm0	���t��Ag�%���UBY�1/��#ГvP��CU�<&��np,��K���r����Nv!����i�\NHh6��*���%��f�d�*6B8���6��&�K��S|}9ZE��No<uEZo�\���t��r6��q��������E`����\�z�YG��"ȫ������"�Ϲ2(Y�ctN�z��t�� �港��$��>��-�>�C�H����~tL�]Χ5��{�����۱�I��i$��	61u*-�> N��v� *)���*��k�B2̄�c����Y6A?`�Kr�Jm�D�|y�4n��[�a�+��k}��q�����H���p�q��3&Axn�݅(�&!�6��A���A��E��Y6p>����R��Q3=(�j�b����]�>�r�J�-
4� k#��Z��}���(k�Y��mt�f?3%��gT�N{�.ͺ���[H�GG$��e��g�b�?` ��>����iQ=�9Kj�����yڟ�G�9Vg�z���఻k�n[���a�I4�5M�kr���s����Ո�T��ۻ
DN�(��c9	%= _&=�Ah�Y��)�� �Ah��ұ�׌{��H�������I������ǭgR�Vi���i6�@ˏ��s/�_�$�PX�<`Q�*_�hbC&�ף�WZ�鯩ӻ1�Q��]ۆ[��k���]j���#ʯ�'�R�X��4h����~�ɧ�R@U13�Պdȗ�Q">�2��2p�MX�ϔ͘��9��N�2�8-n,�J��>H�.+�5�R������&gO=�����⼵R\��c��t�x8��BA��ʄ$�);n��C�����l^')�4�ߖVA�7I+�69dkRT�$����%�q����`f���G:��+/d�)`S���`�h��*7B͚�'���v��4�VEZ8LW��#�h�a��p�ֱ7���&4�^�Y��U+ƞM�28��D�E�ah$�D�s@��#�0#��bHZR�M(�DPg0v������Q[�8�zפޭR!GZ;D{΂;�r�eC��y��0�i0�$���iN`��xU��øE��.�#<���LD�V�ŨJ�ж�rloZdӌ���闏B���rf^���!���6v��\��R���{!k lL$W�B�<ʲ��P����+�qMQ\��x����%f��g��i+�����܍����E
�a+l+�/�#�[��K�XS�V���9��;��o�R�8 s�F~�y�n��<���uج�/c��`�h����K'6��:x���Q�j ��QVy�e�g�+T3�|�o/��A%��	��І-��tc�\7�
����Ks�Se�%q��پ�;u*�<��3Z ܜ�o]�UHR���l��=��$��C4�&�E���Q(�zp�oIyE��?�*avh����l��p�A�F,�P�RG�!�	 /$@$�P�>��U�9q�u���a�@���u�	���P:`�%	�)Ξ�Im�%*�^Xo��[��A���ƀw0	�E�t��W1���E8Ҟ�{r�c
R�����h�/��w�f�A�3������t�D�Hz(� �4}RnI��M���E� �⣑^_�
�:_ic!&�ďd���,^):�G�m��ķ����T%�b��X���,�Z�$��6����:�7~no���ܢMm��0/�b�]��ѱ�9P�~ě<3?����#��IS�y�orG
QK�>��iV���k����܇�Q2epz���}V��a����]��PFP�W/�0�ӼKsQ�C���	07m���i�q�ޫ����>�A���YI���\d���i92|��6�'ʄ���W�`7M��q#�M^yzm��I��$In7#B��
�O @K����Q����n�o�J7�l�e[����{�[!�Q��L�"�S��R��+@��Nsgu�YƱT�˝����DoD<Mgu�Tq��ʙ�I>
V�QG�E2�����W�J�hXr�)<�g_��2f싇��+�??�7��'$�U)g6�X�cʵ���M��@7"��9j��9�0�t;�'��j� ��I��v*D#m_���?�?�]H[b�?=P��Rp䁏d׷E3�A
ap���(���J�ԗ�a��k	<��S�]eeƕف���	��N�ta=��r��v�]Qy{�Wj�j�s?��R^�~��}k��3��O�O��Ed�Y�"�����Q��_G]��I�P i��T�z��*��Ľb>8��Q��N�3�HT�u�}���m~|\)����U�k�Y=z�������ܻ[��P$�*����
��in�}FsMo�P�s�P�� �A�Mp�=��OjH��h2r�(m���`��Ê?z���L��:9����a��ްLuwV�e���Hܓ�G$P�gqO%E�J�𓎅�^]���s8& #��Q��9K��~l�%ei�skj��Ў$�K�I
��)p���W�/h�X�K�p�	�XU���5�XO8�6��Hp�6��JDXA����zư�̚�q��Q%��+5tގ���-���	l��!�.���>�G��ʗU<�J,��X���ŋwa��{��1���L��[p�,��dÏ�
6��?T���W��D}y�.M�/Vx+{�9O�ϊI�睤�;e���� �p�C�C��7�*qg!�}��59���9l�W��7�{��.2�����W�܏��>�RK7l�}S�&~����"��ޯ�S+��nW��?E�{_�[;��G3��'��a����:���2Nvz�729��( *9�R*g$��1��7˃�[55�����
� tc�$=�
��*y�ᦸη0g]�ܙ�qzqf�/�w+Q[e��1Z
ߠ�� �����¶HcK���%��Z�a�9��h�!���P����M90�Z�!�gH���Q|�������&�4U���Bx`�K-�/���qq�|x@���ؗ�y'��@m?��cKō�>�6D�?մ�mi�~wD'[+oh7	�������;�89��ƭ��n���t'G[yKĤ^�Ô$
�����V�3�������L���b��]�V�	;�� ^@��g���4:)M+.}qg�����a؊�o O��E�z�J�����mM���?�����ţgp��ǈ��@�=�ȥ����v�-��%�rOЧIs���V؏��	�z��"00d�`��v����`�y�0M��I"�p��eWy����N6���GqX�C��κ��_�܁�l�r,V�0!�Z�*Y���N,��:�X�\ `;���E��Rw�N�^?��?Q�&\��y��1��kMt�v��x)�w�F��Xn�u���̫���Ꮞt�U-�g�ݤt��+I�d���`�^Dy�9�|϶Y�$d�c-��b9��qT��4ֽzWF��y^fٿ��ÁM`[��l/���V�:w�8�0]s�n��M<���*�^�GԒ,~*��2��K��vZ���[��n�e-
���,?l����O�������i@#!��:O{8iv������1�^�f�]C1�-yS��q_�Ͻ�`��vj�f˄㕴�I�(~-ErB���O�WW<�N�x�~7�ݟ��'��)�6C��1�"|Pbs<G��t�v
,A_���ܦ�
W�).���<��԰ѷ�0h����7�i���}O�zشS�)��Y���es��l_��T�R��M�w7r':i�s0���S��Z�D�=$���R�|ӹ��h�u�������F��cl�`+g�7�ßX��KN�Ś/��? �1�����|�D�%��/�ESF�E�=]\FV������U��}��M�?>������z"�(��?��ɬQ��t4/�|9ue��tZP��t�%�|M�O,tr� ��xII�9�ſ�0�l��YJ���ܪ��Q����<ꍟ%�J��a5�����9,M��]�`�+w��t[%;�Kn�ץ@���xҷ58\��̧���4\��� �:�%�j�9����Y�����=�4iX����pD�ҳ�6�� �1) :{�R��v-���G�R��D�;�ܻpL(�O�a����I2����w�핿�N������tV���g�C�	
���BN�5�p��z��U[M����J��9��
T��Cړ_lU��� �ʽo�b�|c��d�����tz�IJ���TE������x�81
�����ǎmL;��i�/'!�lI��2$U�6:U*15��ho�:s!�-�oD4i|g�������i��|�R�%|@V����û<���a�;>�7#dS����� !`�����<U��4�vԃ����
[.�+s����f��~�"u<���4���^#,+3^�2�g>�U����3�w=ڝz_/��0�}�-���aֻ0���]�"b����l��H
O���V7�O��(Q��2�KGpW��u4?!33���rY�o��[o�J_�V�7Ō;>�&����5��'�{^�H��,�?��)����&p�;є���T�װ�]�YI�'�;+��gs*4��E�� 6��.*K��7x�&��@�mH���t ����Q7�@N� %�&ˀ�Q���C�\��j7�(��Z�-x	!�{x���'�k���m��&��璏�j�*p�O�o'@/�r��z�;o��c�s�Ryq��]	7n����}+���5�U���N�f%�B���z�JTr7�bb�m�1����˜c��s�o�d�Ln���U�����d��VQG���s�F�6�����Kʵ���� D�[T��>K������f�i��K �-P���N����*�a�Q��N�Q������%;j�4w�T�6�C�Bn⃐p&��#N:�g���k�6���,�R��ffL O8����(G6lґq:�01����E:EI�/_C���L���k�X��>�vh&��� �v�+�/:��l��D04��>� H�$5x[73�e�W�J�}�1pF��nNO�d���-���`w7��s�f���w̡�T�Ho���IĬ�wc�9��wI���~Yw��?�Epzټ�t��f����8_��tq�j�g�ņfA�:|���<��sZ�w� �GS%K|�jC���T9����X�`���	���� �}�9b�q�Jf}IH/;H�ք��F����O��(��|w](���N�i���E�s��RL��.o��Q�j���=~fn�%�6uB�]V;T�4�>��z�������R�CC��Y"4(z�Ƈ���p��fd��օ���M�/s��65�*��xЯ�6��� ��nL'��ouoNf+?(~��A����.��P�M��#���#��"z��M�-�Ot�<C���3,������	G.���712�7�l�J*/��!1)���DE� t>��D.��P	���ו}ǁ��I�/�C�h��oJf�#��-�q���ܕ�D"2�q�O�.�+*p�SRk<e]~��'!�F����;0�O0.H�Q��1��t+a~�BI�������,�-"c�3�a���jF����߂��:?�3![j�A��s����U�ʷ��g 京E%PǛ�ly���T֋��e��̞�K�����:��鰶G0-^����� �`�&�m��%�H�1�������-��a	���&��BT_�U2�o�I%��� ܦ��}6,��7"�����`UQ�N��#��f*8����Ze���H	���d�4t�0���R�2f��ù
��7�f7[id'�DN1�D���ҡ0���b��;��7�O�����v�D;Eg$�06�ZI&5$[��(t��A���9qπO��׉�3��� �X�'`I�)�$c8�o�A��.�|��t�	���@���͗�w�`x�y$����.I}!��(�m�*z��b�>�P����ȑ���ڡ�m�X��xv��{sN���E^�-5@��*�Pj�}������C����.�T��i�¯|�D��M�ֿ��	���m����p�+̢�5u���|ڇMvU��	v(C��,����]��Q��	��ӎ	_c���-X�+Q�":��.Lfd;76;IV5��3�X.RȨ;hah�.+KҐg�ƽ4$ �qg'��aj�>�/�e���<�aG�o*����d�z��N��@��R�M�i����'de>��A���sj�.��v�D��'��u%�4�f���{�M��R��V<ȹ�u1����Y�E{K�挪�x�I?eʉ�
c(�T��CNXH�����ã���
�I_����4�t����ɿ]��l��dq��L�V�*&tcn�C�m�xHU�b�
���(����d�X�=�\�<B���<vn�-RK�p��|���ɶK�j��\Cؙ�g=;4�9��,*���-��L�/���a����D���-�=��͡���$69�Ǭ�N�w�2ڍ���I0s��DgE�>l�8Vv���]mf��78��?��	W�>	�	0�,vGF��X�ʜ#�l	y����rߐf"�-pw>��ZA�� sO �ڃr~�����gN�@J�n��]��d޷�4$i���W�HQ^�D �SM&x,������a�'S#%la�!a�ۃ��U.�]����p���ŶSe�2��b/Q(���EŐ�4;����0;ߑ�E�ɏB�@M%��%��:�۱ sa��U <C#��g��K���)� PZW����Rs,v[hd�S�V��T��Dl3��b��y
�ҮK��̞�H}f�؝�%"k{�㋊�Y����C��E��*��C�Тz4�,�fr})�^�ӡ�p;�~��,�4�UZ�1���%݉��(!4�
q�j������~(���b��e�N����b/lH���7;&���g{�`&d�Z	C��1��P4�S�i]5�}�5C��M���T�ӭU|���%��5	�S~zjh��2�E��q|�@n<��O��^M�`��b#r���m��ml��t��X0�4�A*��7�X��s��L�a���C�����l�
����m ���{e*�@M��H�jǱ��|x�c{/p��g��"���Ď��W��zX�TQN!���u�ȼM�+��h�&���d�w©�䮜�G�?�w��]�<���n@�����4�Z��j�v9���ϔ���J���l2����������Gx��_i�%A��D�O�C{W@�k(��|3&�	c����[�!���.ͼoE�~�Q��/���%>�i�_�j���~ 9\���fmv�In��|'c�B�����]bn��Zv�H��Gy�j�5�	�� A��b-�L�*�d�7��^@XP�M�X?�{��t�Wb����z��~�#}�|uL�ע���Xc����@d
g��g�˃����>G��6��J]�Pi����0�a�&g� �[����	.�+t�� �މ��t��\0�);�$[u����?���]�W_�K�[�����r���ŵ-J�)i�4�.z-�KP�|ڋ����S�9�MקGd�h��
��o5���zt�+��
ٶ~Fu���ҷ#��&��g����e7��}�
�m��ZU�{q�x��5�,��M~��\���ҫ	�C�(���p�[�Z#�vä�2�� <y�NT�/��*�V�z&'���;��Co�҄��Y��_`�*�7}��b}0����S����g��g��UA4���êc0�j%(��I���i[���Y�����QpVF-�p��Sc>10���TCx�H\�9s���EH��O|��'_�Nx�������S�`�A�LQ�38D�J?xԄ�Ġl}��k����4� �Lj*�$)R6AY���dH#Ζ���\ߡ�k.n�]�M�R{�[8[�h�8<6v��6�Z
\AH�r8ܝ��P��?���n����5��lV��o�(�O��u�&��ʙV!����N|\���o�#�!�%��r�k�ja�ò��b�`�s�la��8]��\?�I�m���, ך���h��ˬ�;A�$�|S����zXL�T}9r�L�?.�x��w��G�&�:�o�x����D�U�p�n[��s���jw����Sf��.5�6����jB3�y���9�;iG�|��u�`��f�#9��r�lU�h�.ᘃ�A)��b�,�˅�~��9&�WJbd�y.��� ?�10M.d�6�=��A<Q���WS�1
�k���F�UB>��e�{Lg����]��R�H���)!È��"\��ݸ-�v�Rӓ��|&7_H���͆5FS܇k��P���0����Z�j(��,S �g�UC������i�9�`����a$���p�<6r�-䛻�Z�,����﬩���m�4�C1x��Fw�	�T�7�d�= �����|�zw���"I�=L;�~Ⱦ���юm���6,��s��m��`N�8zV�,^|�w�B�(Q����4�A��PG���G���in�&����-"�,�|�i�oQ�v�o|���~�qL�`��1�a�	�cZՙ[7Զ�;:�I6؅�)R3�G��i�I�j�����s)b�+�YPk�ERSv#O.F�<��Ⱦª���z�1��q�� ��{Ns;���:;I�[_��-�?���#�-�M	����ƀؒ��IJs}� (�,�J���D��:ZOA�p��y�9�Ty�z�r?S��8%���J&s�!��T��*�KQ3vp-�>;~2��p�����Qܸڥ�1Z�|?���r���R�M�U��"O"��4��ͧ���ڣ�ۡ��h�����URh�F���T?zh\Q{91Sd����Zb�:N��:�^��2��Lc����4�e��kh�2~.$"^mN�P>�d�Խ �nR�d�t����!ʈ%Y��b@����w�R��{E�YƇ�(M�r����D��{�9���*Gc3	��d�F���.<O�u���6�~�� �O�RJ����*P:/�>��!�ǧ�x=�`�~��`�?�����5�u ���m�!��!�0�Ih�<< �o	|���3K&�^��Q0��-�gn5���^LW��53e�F ��n����̋�۷�p��	��A%[��V��%:�?:Y������zC�?b+�w��. ��y69l����,A�ei�Ǭ���*��x�����cٮ��r� �o� �A�����	3K����=v�Y�*�\ԕ_��Tɽ�0V:Հ;��<*>������!��o��茨���B�#W_���kJ��tr�70�͠Ia,pu�,5��s#��;4-�?��(#��Q&َ��א�0PF��PY�e8�9k�����jĂN%�퇃*��[`}q��E�WV3;z��F���Ȩ� ���8�5�C#�@����d.	W-wu�_2O��;�O9��5PA�W�]�����k�~%w��3C������%�ڌA�5�*Ġ�K�9�ј�n�SW��ؾ)���'�q�O�ν���=����e\?�������mX��Z��%������^��Q��WJԜe����l4[�Em,zN���5~)�Q�
�ab�9�r�:g~|N���4��&�R=�q*_�b<��������f�6�[�"p�Oa'�#���Л�T��ʍl���k���&mŢͺq咃�*T��t�L��a��Tq�{�e����]e?Ӏ��4���0���L�sk��"A�h����0��Ҵ�jz�+z�m}��`84�rKc��xx!LӘa�[B�;��H�\5��'  <��D)�5oZC�c��q∥��w%f�_~>;C�f8��ӣ�a��YD�(��$`�É
"$�v4��L�0�P�↰�˃�m*���<'D��{	`%�����H�l͂$���\R����!^�s��aqYᗠ0N7Q��0I�� @>O�eW�d+u��K�-���Pk,ҏ3�g@ؤ�ʢ謚/k�S��DH��ҴZ�D���F��'�6� ��O1p�_��U! +���%C��|�,���j4Kk�̧CȎ�էAЫ��4Q.�͡�j�b�S��5%��XZ���R��`�*z��MTJѯ䈢)�l@�Q�e�{~��*��~�������z����"�>,�'��̿Uu��������Y�I�V��P,��ޑ�7��z�4MXpCm��)a���BJ��NձR���a��p$Q�O!֘@����)	KV$v�c�eJ#hԒK��_jugw=�K�|<L��_
s !;���H3q�� HЮ:��%|_ؾr{��wU��\��CFF$��ϖ���yc�V�(���#��W�
,��)��橓�R�K��餌�NR�t��YU��ݼo�?X�'Ez�>s;��N�����iƸ*��>'��@��s��@�W���8�?�����t�󷈍L����r:� 4�敾;�Kl��J�������P�,q����<7�?ڡ�q��Z�����ù#G.�nF�<����\)D��)�LV�n=ư���D����Gb�𙊪飲&��U��d��eȬ������ w����M�����c��}�I�B��r}L�*���is�q���v|)�[�y3;B�tD�תS]�g��Yo?G�L��k��~ ��֛>��"F��0 f�)1	�;��&��n���Ɩ���JUdϑ!�h�2��ˡS/��$��X�+��\�l�I�rj���I�S��r�j"�Y��y��(���'=ȔN�=��ߪ��c�"Ӏz��b�����&��p��� '_�~ͼ�=�6\���٢&Xg��H"��ɟ�,�����:���t~���r�
��)F`4o�
ϘM��#_6��V��ww�+��C/$y�����%5ƹ�����͝=�L�ko�g��r:�<�Q�h1�D�?Q�2�����+���}��|ݞ��n+�𜈆-L�y�871�]�[�Jǻ�F�C�p�����4�*�|���p��&u�]�C��ў]��zQ�4��gu�"to���$�Rҳͬ�F�ʥecF�v:45B
��{�]r�h�(��sQތB��q<\ڔۿ�<XuN���ܬb��O%�"���Xǔn.Ƕ�#Z�������M=�wNemY�İ�?~^�;]�.��`�Di>�J|4�Zuc8�����L��jrYk���{���]J�R����B1�4�dQ������f�GwRO(����;'S�����o�)of��:����hcG-���)�%.������y��\�\0	�b����@��qS��b\f�e2��*�І$t���H_�'���Rm��,t1��|�M�w�F2�C�y�34��a���Oýeꉫ�$��7�[f�5T,����6,	"��ˋ��r�D�䡻�Hx����&���Na���o���!�M�tX7��ǫ�����n2-k;�q�<�R�q��w~��#.�\hRiB=x�;�1�<V[�}�X�VƵ�_�IXxV�Ƈ�B)gE������M�4�;���^�
���NZW��T"�{� �/lw�E%��G�.�S �LϺtctz|�n>TF
�D������MϙԖH쯈G�?g��W�q���~Pj��#���	\ퟜM��nO�g�里��)
�H{���Y*�n����2]e ��<�n*X�������2b�b�~$V�+��m+��|A��� �?�-�,���oq�<����$������\����<�6����	h�D�Z��x�H�vp��~ؾo���I�	EF�Ɉ&-��ѠGǆbA4���
L�/mN��A�c�>��g���;�l�ϕU��;�"a*�=�c�ˁ����������$��@�����y��~f�|����̈́`�R�x��V&�Z�q�r
��_5<W6��=���<���˙�<�R�#5��)o�<"#�Ԟyˢ��m�᝕�	�.�тX��ۄ�G�'��Yۮ���gfÎ��KS�?Ȇ��[��8u��PD�?��ʠ�	ٓ6����S; ��Q"�����t}+m,���S1��������|j�D:�b%#�j�b�;���g2v��ɸy܊)_�@G��&�6`�słz���X�m�p�~��JS�5��C�T<x���ؿ^�F���ܱ,��T�h�K�VR5� X0�l������e�ATuC��*n��x4�L'&���-�B}���l�����67���ߢ��꬯ T��E	�l��ՠf��Z�V�/3o~�od6�N�4Ni�e��-z��Gh�D�R�ß~羟(����d頮��t�4�3�=��<@dy*Fu���^w��b���#mǘ�[Β�މ��p[0#�*
�`�On4��s1N:jgb�sϊ�
����Я�)>Dx�|��|f�aN�2��GēN'�I�{T�1�8 ,)�i��R4@}5Kh]e�3�_BP66m��!a8D�'aS#�u�[f�RF3��u���6�6t��̣�˸=b�dk8s�A��-}�X&�?�wQ!�i-�?|8"��������j]���:{D�F�������� ��<���� 2t�d���9`�	}�Y0���P�k��C���mm�JS.���Nk96��tan��f���;k��_ʡ6�D�?�Nf����+��c5��z��kfY�)���X$�~x��H�L�\]�L�KG����{_
E��[�8����*�2e|���u��9���
7�}F��OM<��6-��!gy&����ǐ��@-���JVHK
��b��ݟ��jp�<���A3���ͧ�CG�q�Z�Z~Z�:х[�&:���:5��mǅ$%(G�Ч���փx��`/�����������#X�D��l�ϑ���k1N�{zX��
%i�E�ݶ��h�gz�+��N���^Y�L�������xl�07�����*�T|��o�`�Tr�J)\�Z�5��������Ͱ�A}��U�)��ՙ��;����0ʿ���B~,�BqEŅx��Ę�o�4M�#�i~2��s��,�C������$v���@���}GF���"�J���y�M00L� HO�!%5����qz��n1�G�Ⱥ3�:�֓��Z�q,�L�����2ʸtnI2<����H���hF.����L���DϜ�WX����IA��yÊH}|���y/U���Z�Nh��94����8N��7?�tR�Z�/k��@�_�n�g94�W]X2D����3tft�V-�����ٱZ�&�o�(�B,ԟ����]��2�ټu��N��A��N6�_���W\a��(k�����~<[֔�ļ�>���ji=���tk�/L�.���������=��5�9p	q�)�$�7K�\;�؜�v��!?�����1i��
Im�I��D���T>���
Db�#T��0����x�]��LO��ܪDJ^����"/.�z�΄�8��w�����;ek�G�G��� _��[L�bt�sٸ
r�$ʄ����,���)3ձ��;��3V��F�a��(�&�ۣ2���yGQ����JIz�V�Z޶CB����Sa�0��-`<�S���\#
ۇ�[M��1P��י[�*^͢�UU��}���-�b� \��wQ��X�a�q4�,�f-�S����ȳ��eq��5�ū�F{V�GX�z�Zv�4����G�^T��x&vPz;��ak��)��H���D龶�I%�A,C�)��G��Ok���X�]!Ӭ�`�f�V�,���ִ�MQe%�-|�3)�#s��!��b�c�V6��0Tw����#��å9)0F�A{J8y�AC��i��u�16uj��t�%�=���������P�s���PL��En��Y�{y�6�O�I�I;u���E���6r9T��(^�$3v�����4�Uw�?'�r���.�<"Q�KD�gKD��	ݭÇ�e��:BE�3����ֵ6�a���E�N ��P�"���2+.���ȫV$Ɓo��NP牋0q�b�F'����;�.�T��lxH�M�4;���'�;I�DS2��,(RY��T;9����q7@��-\���-��Y��.c+N`8����ȥM��O�R�tv���w���W��V�WS���h���=b)ׅ����g6�+���J���"�W.�P��Y���vkZ�=��Q.��r���-j/A�������;�H���S��t��<�i�V*�[�@"6��M\ӂ.��/[,?�"��h�;���Bn�&4�w�y����"��k�:�ӱ�ظT��D��QEWj�H痂HJ%#fP$��Ŝ5� �%c-2H�*8k���������B��"&ՙU�A	u�s	�$�T���a��+��nW���D*#U�%ˋ��T|!Ѭw<�s�G��Moމ�Ϝ�+�ٓ;����u���5У`f�#��� ��'��e�)��aT
�г��FT�`�y}a�J	��A�����L����wJ�yi?�Y�Ԛb� �s�������,l&,�i_�V��"$�K���f��/��͡)����,�J?�Ʒ	{\�k/N����w�o�� @�~�e�V��K�����V���Q�8b�8�-�G��J�⥘��u�-4�#]r�n�����z�}������,<@-�jT�NZO`�U|��w ����K��I���a���wg�e��u������0n�D8|�G��CVL��w�k�Y�ȣ=��G�cP��ڪJߚv�Y�S*Q��T�5�vy�D�"E-x����m�-��C�3Mn�,��hS��m�*~ӻ֚1���#h��U�)z@!"�
�>���UTB[���i�stJ�9p��W��]B:�G-�$��E�y{���K5�=�����:`�˸�ޱ�K��L�}_g�rfb&���8�{?=࿿�~��c�҇D�Ě�B���P�=��MN�i@�>�г��Jn�v=�u�uV`�$�.���O|�{�F
60=��� �+'��_�eZԙ7��B�Ҿ�� ��tS�0/��_v�����d&s�<��O���F��$G�W&>�'-�A.DmA�K�5ё����E8)WE�|���#^���ѡ��QNMa�S�]�cx�����<9msI�{h�G�n1"tA>�u�5��s��+T�N��'��8S���K[�x1͇�f�Tl͂BD]sn��Y�"d �NW�HKg2 �����PC��z��5���������J2�W�,.]��<<��|T6�'%�#_�6_����+����ӱ�)Vd�u��O��cy�7��� �k�m�4���,�k�P�K+� Ɉ�w�{C�Vyc�5��o҃"1�:�p��i��F��q�D�0Ȼ�2�k,H|T���,�j	k�V�WA<��ƢJ%����;5:/��WwF�
�A�G�`��գO酨�!��:
v��;���=g+:�=*�O=Ql�v��r��s6�9�V�`��B�r.��a)ify�G����y��R��*+��@�k?��J[�(2H����B�)���q(A:�xiEF��s��|�mu��U��@�Xz��2��ٱ��z���(��@��ꔬ:�y`T��k
�q��r�?2�8 �)љ~@0�M
�'V:Bi"B;٥c#1<ǝ�я2�*^i_�#���[��ֱR�嫈:߆b�7F�jT�b���:f�uop�sGF����~�$ta���l? A�?��o^�y�����C�t�O�l�	F]�
DLJQ`����VBw�Xq�@���#��� LݟO&l�a�����d�ô��,
�,�2�uJÓ�.�F��^� �^%IT�U��}���չ>@��5��-2
KP�،}�kZnp�l()Gav�LL�����Z䚟 X.%��q�]T7�(5�Q&��"��ԖA��Q�H���Z\)�&_i+s���aN ��j~�}L.�n�f�igm�aI_�)�Pp�x�i��n�2�d�FO���@��L��h'f��8��Y��!S�쵠Z�&aɵ��7)�66��Vi-������Fنy{��w�\Q17/�HH�֣�Pg�Ј�>b��a��RK�Ea����,Xpɲ+��kyu�(�^��!~z}��+>�Ī�IN��**�{\áf}gv<�!"�-F��J�;B��Yo(�% }�Yv-`N�Gzʵ\ܡ�;׀|�KwΚ�^#&}�\�q筞�\���`&����Q]��ָ�ow���\O�n"��^��Oyf��?����a�Dmږ�JEQ���#�3ص��<�|����n�W߱�y8g�����+�{s��H�FN��sj�����Y��It��Ђ�?ҵ��Ƣ��#%w�����"D|��V� ����a��OO����c��~G�%�u[/	r�P�;��픯��gn_�É�OC�AGL��)K����'�U�a��T��܂���7��B�$��j�=��;�j�jA�Z��|+v�o\̲/��蓁M���8��6[;2�%�\U���m�dr��d��O8��F�x�~��b���^��Z�3�26>4`����� ?#`��i��^�H�~��N6��� ��ȡT��GPU0���S�j���N�j�0Q�0�2<'�=��E��w�	a�p��f(������.��	���3�2xd�,���?25�T��X>\r�U
��FW�&��r���76�:8�~�4k�/	���(0$2kq�y]{pT w:��.DaL{.������Ftxm٧�V�2�$�>⅝ӝ)�k���ax
�m�ᑐ<�%���+�&�jm8��xn���=�����O�}�H�M9@�����ז�l)�~Z�޿|?�.\�����KE;��̰_�L��(4�n�so��R?g�g<=,�'(�s+�S���F cy_֭�Dm���d�(T��G�q��*~j�R�f��wN��� �O����a ��qۡ5N�e��jJ�� ��F���Z<O�Kb��*4?K��F9GR����orG�F0����f
���LA֞t��^�ib�!���(�����k���u�w��EҐ��wv��6�Q�"f�7�IW/��U�54L�l��B�"�mR���Y�%ONQ\�|k� ��0��wB씭��
��)��Uw�y�{F�D�MR�q��J�	��g��33�#/��[v2�&p���tmy�b�U�n1�7t0�{�amH�SM�:D��ڻ1�OR��D�
�**��Q��J&?�%G���,�X�6�fk1ڱ�<�?��N�P):�5�p�A�V�< Kӝ���]��96&9>b)6��/��7FAR�� aR]h*2U���?L�<D��UAI�\���0���7n{�]�"�`��X��{e�zM'4|�ȿ��5���@�V'��ߒu��7����G�������X��v�h�#L߲c�:�~��C<�[����x��R����i�U*�"�Uג��+�!Y��F:ؾٽ�������-11�&�W:�~�?Ȟ
�RX~U�����n<���	w����0�kw׌S[@��链�rQp�����TM����ll��h�@��
�Uc-l���W�/c"Kq��yL�p���aH{  az�� nu6�����.8�'��L�9<��fߡ�q5���/9�S�*�R�W+�� �o��Z��\��v�R��"�՘ v*�Jn�5�����c�[�L�?"�@&�ǲ����e��.�%Ä<�6��=�軪��wd>P5��-b����X0�	��R��ld
�gۡ�;@�zͭp*�����������N�����W�� �"��ㄐ�M8z�)�`�<H���SW��u��E���Ӊs�E�-�c �I�	]���ŕ&;�o�Q~O\�1?�N��Tm̃�Y�5�	Q|�|O��zz?��h��3����|�~��#=#.��^�U�
��B��\G&��G�ȭټ�TAF��m��@����Vm����_ݢ�:�I�i	t���*7��	���7�`�,m�sm>w�5��F��J�4��ܵD�iU��ޫ�i��c<�����#. ���NI�x��ia&�&kpT��S5[-�{�����2��dE<�va�;�Z�����zUK{���<`�i<�A�G��u�+V� ��#I��=pR���X�z.�5�@DpCt,P��k|����J���(K�F����{���)�t��0��	�F�y y޵N&W�_n��P(�;�c�(��ڄA��IK���&w���%�c5%9ڶ�x�(َ>��l�j��"gU'��}���&��q�'�:?)B%0h���g��G�l:	�s�a�#�+��\:�	��6"���:�8a��[R���Z�lw�6��inPt0�M���h�<��:Lh�m�C��_��,���%S�}
3��%�.������,Y���X�o�[��LM'��0j(]��N����
��܁ B³�3{� ��Z�S/��'ky�^�и��?�.�n�;��	���e�����Ѓ�i�%��Fɹ-'������Z�����j�D��q��l�-o�1 �dY�Ԝ
����h��k\^ސ����c�5Rږ���a�7EB� M�k�X��>�Lk`�ē�EC�L$����־ǒ_��;�w���?�î�����������+� ��Л��.��ﷁ+�o\X��j�!|H�E��u#�6@N1�u7Ȼ2�u.�;������O:{+=S���h�U��@�4�b�
�7[��H�G]�7�s�����x=�����d����sdi}��|^��eg�
�-c��+�1(�'�yNY+ٜ�y�(��qΔ��̗_���?g&�`["u�	���Z�5��h�~��9��&ˋ�=.�lê��B
�q(����z(,$(OT�KE=�]3�r����<���I��F6�4�ͽ]�P)����I �#YO��!�L����u���?�Ss��Q"n߉XŰc\�Mt�cX �5��hHR�b�(7l�)�g��X�� 8i~uu.�I�j�!�ӧ��^?�o"�Ú��Mn/?L
�)��5��Iv��lyk!��#�Q�N�[���O� ��3��
�㠔i��ـ�@m�%[��΀�ɻ���X�q��T�7�;c��WR��4n������ERG͊BF��N/��t|��A�nlO�����/k�x�Ø�/�0�cf<5Z	�Q<��;9ry{K��:��i�/`�&��w@�Bi�M7�*ҵ:��I7����{�[���Y�ێ��P�;�V� j�[�*qM�� ��L�������Yn��PzI�E�ב�I������kV��v���}K�Y �������T_6��kqI�ue�i����T�" ��6��qwս���?�����l��ث�EJ���Bw����y�ݯ�#X��袄�<���D��\i��)� �����Tٲ���$��7R�}{����b+�MGW�B���!2��	9Ce��ɂ2��ڒX�D�'�;��a�K��V�&4(�Н�Z6�-�ܜ�8�
�F@��_���Er����������Oε�Mʘۉ�p��@�.a�����d�#!¢���Kᐐ�w����0�N�)�ϛj��M���L!��f�:��ү��_�������N��b��4�?�ݍ
���^ȏ�V�E逸9Wkħ�Z���Da�o��j�ֶ��<���-�>FR���yz,G��VY���"5���Pթ$�,{�t�M+�s�J�s��[.��c/.�'-� �F�|H@�0�����M���;3��3����W�bC�kC V��Oеs���|�w��)Y���K��ct��³��c��@I`�yG�.F:�4;\�<|�[��l��&Y�Іo���VL�W�z'�����d'_��V�/��;xr{*���x�n�U�3�@kX��7K%�cI�똡GE�w�������@�v�PPP0f�%��P~t[��U"x�d}]�/��o倎���oZi�-o��R���P�i@+!`�I�xh8�s��_��)8$��{>OG��Ŕ쪐q�t�v����k�&��������PyZ�Ty���d�U3"���ZHrQ6m�sVjw�,t0��j.ޢ�B�?A�
�4LyJU���#���I���{�5�B|�	?�
�p^��ےx��۽8tR!xJ�_|ŋ|d�fXY%���!gt΀��)�ɐ��};�<���]��N� {�����H�^jU�w��� �&ÞI�,����sQ����W�
�a+��������������c�"z-�����w��0�
�����w�7���l�B��YX�m�m���[0��TۨI� �ꏗ��}qr�F�X��C������;+E��x�z��݉�ߔȻ}��)�f;��jQE^�Q(�&��-v(����z�hۙyZ���I�,��]CyC�;n-����B�Z��?�e��~y�J�Df�t�MSモ�u����.;�P+�Q�j��|m��M�V׍�d�OE)�	̤H�"�ɥ��}4f~aiE�^0]x$�}��I�G}��5m�>��ٷS�3π��)�>��h_[�>����](̊���R^�V���>�	ߍ�}���#������*�:��^ &*�=`^yE�Eۊ�9V�7՝b�e�hj. .K Ҫ���z!]�j�_]����_t���Q�Se��bʺ�|G��[t�;�Y�qv�J��ǌn�>}�!p��2���?�kt���sE	呏�	%aR����3��-�ΰ�$*'�E���T[��p#��Z�}Ӊծ� '���� ��yA��Rk0�!���|�Mț]<�g\s��g�A,V#R��,��]�9Y�Ku-9O$�q�����hDh�,vx>Jx��&t���o�{=Z>:�ճ����~��7�8��3��J��
�����6�)�R����37�}�v/�˝�*�=N�v+�Gǆf�%���H��P����6zSd��@�S�-���Qh��D����d� e���v�|���s�f��>�F̫���N�)0}C�%$ҝ�s�o����i>�>EͿdA���h��%�㗏g�q�|\�:^���v�y�'�R��a���8J#��������5<���TEY�vCr�{˗WG�RI���U��>?�o�!�	#���Dl��&&�uS�Y~��M��7$b���;��鰍�H8^�Lm�`��G���5��$;>��6u��FU��g�	�����-Co��g��߂��b��ͨՋ-Xi�͗���%T��뼑ٽ��u��x�t��kʱU:a�^��\�<Ylo�k_�_�H<8��n5������KD���\Y�;�@�e@5Z��7	r�/�ԧ
�;�[���3]��B])��'X�P�+�ܡ�&�w?8��_�3��������+�����l�
�i�3����s��נ��]��/z8t��?�����.����Uزcg.��R؃NH�ޓ����F��0�!��/X�V>�����[��[�x��u%�E� l�����3�21r�	ZY&�[����K�1��q3t ��=et�c���� \/S�9�E��þ���}����G��CƐ�?kT��~��>Q��s9�{�ˊ�`Ͱ��`��G���g�J�{45>g��{q�怕f���pLp�?J�SxQ_�~�� k�/�b,ܬ�H�?�y�@�T�4�:RTdV�e��fT��/Gt�B��
�2�Ŭ-a�a,l]lx�B�=�����?�IC�(�U`�>�`��ϖ����x���E�%
�w�	K�	��(�v���࣏�5���b"������f�1!M<TM�X,7��+O�%黆��W�p=�נ[�)� ��Շ"�b��,��'�<�r� ���È�~��pC�ރH�n���|WŴ^�
����5��y�Y�8�����>�GnK���.tf����A�k������#8�X�SyHZ�d�o�����8�)o��A��O}f ϩeVq��ݝ00n��bz+ �5Sw�4����7��0�\5�:G�jڈ�������'NUL�٧��p�խ�`���_���:�ZPM�1�����2dzQ�熦�H���-.x�#�7�ci0B՘�v��n�#R��^�Ⱶ΍g�
��؜q��,��%%!���P�	ܒ�Z���!�������QK�j]�z��QBX���UJ�Xoq��5~�����~�ٛ9eܓ�ZrU�����1��b�]�|��*���y9�����<۩�0���-SU�$- C#��Bz��/�8y{�~Kk���H}��.�q��gr��Rnd�	F�K�PY��o��+����������r?���h ���� 
e��s���V��גi�p�1���8�S��Fć]
�ѳ.F���R{��UP+n�����������3�h{ve8yӔ�.1���$�o/�
�����z#��E�8n�[��V��:HR��8���kL9icp���
\��UT��X�~Ȏjl�<ʐ7޾��PW�N�.��/�S�2�k���mc���5"���̾8݋�G�!���W��ec�
�/���m��D;2�&h�0��,zq����^eu�gj�d&�0ч.?/���k��Ul��)l��y�Vyk �.����F3�^���g-;=:�U�o�xϞ�'�Mܩ��Ơ�S���k�L���~�^g�h ��)��� �Κ�W�e#c1p��x�I{�/�1S.�]�P�a���H�X<1�M�P@v\D4� 1�y�^���;
oR�|�-ght���a�
{�,ކ���	�g!�z����^>�^��[�+w�k����wƐU�^؎��'"�S<�7ES�@���,�.�M3+�vI����Ax-���^�m�ǁ�b'���4�E�0/��N���ݼ�m���%c����?�B_p��P(�� r�ux�t�����4�G6L��M�@ <��&��|�~���D���S���WT��;#,ɷ|<��(�T��;޿��h�vfv�OzW�r�A����ee��t4@�]-j��8�L�tǧ�Q�ޯr�].�هK���C�Ĩ����lX��m���\��+9����D�W��o�s]����WP������1h���Ѯ���k���?r����}�g';��WeMn���} �ka�U�����+$���Mوa@�h4��𝭰U N�y?q�e.���r��N��j촯��"fTM�.�4cX<*���\"}pͷ�E��@@����
_f���M��Fq�`�
@��?x���� ����5��1C�h��t�^f���&���E<$���[ʍ?'��q�A$�v���5_�Z�ZAE�M:�8^ �@Q݅����"��lO<7mo���M� 5`�,���$�~ő8]�{�o��,��Љ0�p8oV?{[z����p�s�(j�dKL.QЬ(r�X=��VL��t����,4Ă���Gc��9�4���`��l�/�iN;}�M��߷T��7���T�݆"��P��� ���zm�Z=����3x�M���vD�߂�����ن�1�X�1��J����A�֯��,�&.��֪5��~6(��M-��\�� �U�;�u�e�8ߞ uNc����Z�������g�4!� T�׻�p���m�|k%�Ʒ�?1�q�ziFT�ij	�U�ǆ�v5�.���$>��k�/�Й�AM�A��#�Y�����!��\�Em#��Je�Ti�*����{�����Mq�LO�
V��)!��^�l���!i��!sS`)�X[������k�%�dM|3��ڙ�[M&���k�u�":��pD�M5��t}>���nF��8�|,�9�����(�������;[i!
���C�{��D&��]e��#�)~֏QȈ�j�EH�P"Jrf2d��ݵ��G�H �|x޳U��=�f��Mz6�户�:�`�ZP���M������=d��L:Z��/mIq̸�F��Z^���f�e�i�yS��Z4OFa
��i(O! �@��:��ķ���i�W������7q��C�I�Ƹ��e�;t�jD�Bw;�t��۟g��:�"$/�C��
B@���0G����FyU!=]�z
�[�NL�
��X��$��Q�`���`>������̓Kֽ@��g�P��"C�ە�'���9���5"vo���)� �16L&Ic4�4��1]6��n��� 9Ƽy�#����ux�1�l�-��PƆc����> �;��M.�J�A�F��a2u��i���9{��|��;|�
 Lt*N�~h�U�B��������f2G�'��VK�9S5*��Fہ�FHLw��i[p��ji��mwc�V��e޹ڣ�&t,�d�� #�W�@W�*r]� e��&���̙��b�g�'�l�B�6�L��a�8�5�{4qm���} r�J�nc-�a_����E�p�<�y�U}�K)�)��[���@?G��Zv/�Y��-�3]���!��X�T��b#�4���扷OS��R����RԘ�E�脉C�����#,T7h��8ן��4��׀�����J�}\<�$����P�I��oIh�_�|�E!QZ\���$&8y*�[����/��F;����NA�:���'H��qQ���Ji�
�a���.\��N��{����ݢڄ��_��@ƙ�<A�vǓX��|�����Fc���P���\$� ��Rk����pB���
75Llo�=1�۰O8}U��f�Y�<ӷ;G��"���,
�B<j߹)�_3|�낓�[љ������1��l.f�����'�9�;?�VQ��o��6S-س�燵�5h�iP�<��2�T+c�@Q�2~�����R�`�uUw�����|�~I�������XBL{,��ӭ.;0��'l'E���6a��BX/2WM��v ��jy�x�E>�x	(��wƃ��Ĝ��$�k+�4���3�t�ڋ���|KJū�
ٱѨ扟5�@2$T�,sX2��]��U��{�5���'\[�$�]#"&��_�.�����ߴ%� t�
�Se�iL/�C2�^x��|P��s��e<��I�8���ȵ}�D�Sx�L��ڥ|�Y�FC]/�� �:r�B��pW���DD�V�.��׏c��qq3�/�T� �%�� ʙxmGsA����ݴS���lJ�#Z�'I�<�(;s�h?`b��i%��D\*��z1	���<Rٕ���!d�5��1ᔑ��b6�|���4@d?���`����(���Y����}�Z�?r�a�1�,m,��XGX�pds^�P߈��.@0'�������:�ȥ�>�a�ۦ̈́�B����H�Z8X�.+݈>���=��"�S��bP�P��\j�%��к>aS����)x�*����)QuG\�QA17(ߘ���&�%L�����Y\�
���f-j�7!�����ί(���/F��qB)8���3*~K=���
���O!���q8Q�^��	mK���E��
e{�i�|�+�����q�S��ݚ-�����ĔN����E�s<��
�1��%7�cs�J~���W�% ��@���:�����Y�,���~md'_���h7A�Ϊ�)���|8~ z�	�DN�UT���q�ρ{9s.�G=�ǘ�"3�˛����⋉l�2�����Nw�ڀ�0��nN~�Y���-�)n0/f�u5B�]�T�aHeѴF�d��ҋ?��eO�:�ps�������X�a�t8��s�ѿ��	�ځlf{���$��k��WK8�&tQ�g,����a��ɹ}���v��<i62;X��w}�O[��Z%����LZV��j��O��a��<K���1.�p�T�c�/�V+a���� l���1,�׏"��$�8\��7<�b�:�rE[���:��jh"a ������3�i�� ��+
�/�RH'xx����R)�6 E��Z�(�Q̯�&p�^BC�`���p�R�$�4^�����6N/0y���x�C \_N�疅�T�>�F";]�8�+��+�2�d��R$�Л��HQ7�	�;���'ǣ���J���Ek.R��2��<dI�-l���4����r}����ٱ<^��]����β4��h֥��[Wh�'5:�i`�ҵ�����N�g�a%�*N�ׁw�P�wX�*c��K����`,��ao��ѡ`���*�aN�R/B��NY��dqN���L��7c���\��]"������u$<�1���d+_h��邒�s�������$�]�\L͚�)��^eo�������� 5~K�Jg0� δ�y����@C����v��I-�[V4K���$?I�l��d�t��u�׽����/�?գ_��I8F�9F�������F<E��]�Z����\Kqq�ݑ]Y ��G/�}"w��(%I��K\
�`p����r-��!����P73�x�ρ(v'���r�X^���{�~�z9��x;Wd-�sP�#��	�rv<8��W)���62�x����v?�*��v��)�!FE6[i��H�KE��4v�t/�%��4Ў�	gmw��}Sd�����x�/�$�,�s�qE>x��3�H|W�}Z0�I��G������t˙@5�R2�70��ȴ]�8��N1'Y+�S����	߮�\���r�qg���C����L��y�hT)bEA!�C��6���L���	Z�x�R�����{���i���/,�
�*��j甐m��凧ҳ�+[��*n�պ��{�kD�6�.���L����2���s�.��2��]!1@Ua��e����n䛋\y9�a{�l������޻��L?�
B�_i ��M�A?��m>v�N<�g�{V�s���(~F~�.N�6��I����5�ɭ��Xvb9��1�{����>�%l��B,#.��9ƃ_�#[�����roK������b�G���'�4�}��6ב���W�;�>�;ܴKϱ�F�g��e=:���^�2�z΍&&Cx]��:�S��ֲ�����#��0�`�爀���y�&Tp���CC�C&��4�o��L���/~i��Ի�t���u0���S�o*
6h)�yG7ri`�"0TG?��e�6*{A��A��'"�0����M%PbWv��I����>6�����32$r��;����9���K�|=0"g�eA�m�JeIhPaFɛ��j9t7��@�#�J�00��o
�	�azn9��]8��?���c�A2,��3nyP�o����N@\8��ig��$Y��|�/s�1���A��^YM�\��,����5��ٰ�=�����s�0.]L���x�qkJ�<`��=�#��S�-�5O��Q̒�F[����o��ʧ,K)�W7�(1�����3�ʾ:!��+�ʬ��Ma�"���R�1�	����ܞ���Q�O4���s�O�����E�@�N�)_���H�ұ�2�*���&���ȴ��s������:À�C*�wrc�Iv���O�,�@čM�0���o�,��<�̠� �[+Ud�OL^ͨ���c{���w����s󦈃�[~[�D����6�����lg��G.;�Xpܸ���[��xRdL|r%ە���o?dM�����꟪[����	� �4�-�'{��/<��; ���}0<�c�G^��>�]M��Q;(������5�K��z�ɯ��]P�_�����dN= ǚ���b�t��i���6��W$u��h'��v ,��x�Oqk��D�ӖguѴp�-�t��m3d�4(�l7����,���pVf�%�_��^vϮ��!z�3M��F�50��V� ��(R)X��j�陛�s�/��IEn!���Yh�JI8��Db'������:������4�؜����\��H�\��_(`Z��D�_ͩ,>O}���ж���c�����pa�Ie2�q2I�:=�B��V'�F�}��1��:��Dal\j��!� ?�o�(��<�'ue�`��IZ�F2�v�9 �"���?�����i�~7�o��wD�ǐ��ZDe@�E�RD�v�o!������P�t'�3wu�b/��kU���>?h�EI����i��@�!:��7\Ew<p��%X�3��1VBP$N~y�$��I79μ�!D�o�Aκ�.(�u�)�HN�1'�>�A�y'�h�,K4=}���GR19�̆��G���T�ՋV�/,�%_�A@a�N�" �	d�#��k�vT�?�YS[t��'�I�,��K���$OzL���p��y~Z�p����m�^!�຺��ـb�[��_�r�Pqn&O�Sc�4��CѠ�7~�:Y�Ԝ��@�0�FͶ���WR m��PhӤɧ�?@��%��� �(�O{"���$�+��8�1�W��e �G� ����
?���n�i{�,�{����*��&G��`��{�����τ�	>�)�83Ok��5c��3uX���g��#�/bE�@6�I[ Oح8T�Ȓ�'0I���1�,9<��KBG�	�s&R��V/�J��)]dJ����p���\6����l�z�Q@/�b��9ٟ�YR��e�ڪ��p���(ߍ ����z�v��4Ɲz�%?ƶjsf�?{E��p�qJ�����m-�&�Z��sB[�ޚ�pMX�5=q4zenYq�L�.��Hy�D�l��${���!��0�����%��ZHғPt��@�X\�s3I㪷�=��AȦ�?�l\��G�Bm��	 �1��δ\�4%�����x)D����@hܻ��ݝE�3�=F�g�������͔�sC��F7zx;��M�t�|5˅��fز��w ��Y�6Y�q^
�	@v��o��~Lo5�rncŶı=�5��W��?	�����^�t*1��"��.c�.�jK`H��`� Jw�AU�Н�e��Q=�a2��[W(��k�_���МV�q:[�������v?@pϐڠ��YԽ8�)��{!�3�f\c(�>�^�ƃ�{�=����+���R���3
���i��x�M�K`@H����,�ʲM�z�u_P���g}����U����æ�� �8<�JA��S���t�(��('���$e�(%/�W�v)��'��u�h��+�������D����vwv��nx~�P�(��[[��;S�ؗ�d���V1�������0D�쇋X~�憶ң��b���#�yV��z͖dD�$)ؼ̍t:�����l��w*s�V�`�/�o;M���-�+S���IE}~"dͨ"�������V4�}�wC�]��?���nƨ��|�-9����,c)��g�a��8/]T�������
����a+�3y��dz�\�} ����FC�ػO6��D�%�s :�L�t�ng�*�D�Aݳ�gk�������*�
���;<ǚ�zo鬂t��;T�N���!=!��rbI�h2�n��L_��Y�w�Ɏ�g���t�[�/�P�Y� ���ۘ��҃���D��z���$�|��5n�i�l���Vbd�"�{�dx¯���F�� ���E�i�����IM51�@�a�� ����p�f��|R"�~]��W���0��> p��-��U}�ެWfJ=����å�P�k�~���3�¿Δ�;fV�	�T�eѐp�Zi��:�/��o���ܩ?sj�"g�Yq�O0t\���H]7�÷�Y
����o~3��T(�Ҵ��r{�d-���7�7w�� [�eQ�������%v�Pa���Bi�g�b�Z]bH%%j�r��2^x�y:w�X�-Ɇ��F��}�ٯK�	���Q�S��gA�	��]���|hN=�ڧ��;9�-H�׫��a�z��/ Ђ�e�r~~��d�
l<g<r���;r;�)�l�_��ެ�eD�Rfe��{�H�+��}��1��;�g%ч��ζ�����< �_3��F~�Y%�	�A��2{��Nz "��9�|b��s9�9z���$�p0Bj*F�Qu��/M`�{��A7���������m�\c� þ���un�b����߱��ըE��O�1`q�yO���i>���5$�L���P9��%��q9�f;�%�-��A-=�1�'��H�͌G�ّ�l�h�OnR��«�I�w՚� z�֛��fp���`i��E sL��
�v#�՞��~@��ם�k`-1���B�Vx�Ik��_%1�M��W��]��K���[9�Ǫ={	��� K��A�Y�7�	�Ր�)
����(�[�6�Df��hl$]
��>l�j�W��]��?)$s��&㭸&�'ESF�P�ޡu����Y"̗�������Wb�/�S�1s��pC�F���J�b�g�]bSy`'����K��Gǌ�w�m������=8�r�O�Ǧ3A�X�p��I45�>����J�/������ЅL�V����!�k$;>ؠ�`tz�7A�z�6�6������ɛ�Q IU��ǂ���]K�P��
�璤^.`�U쮍鷃�Y�t���vrs�>߸��[4#����r�-���Y�u��A?�Ρq�{�O�z�Md��)e�Z� �&�D���W^U4��ssN~M~��<bkqgn�����mi@�����u�.t[�������L%XM�e���j�1����,��m���q�J$��:/k51�"&�2!%k>�@4�13�:m�f[�!Ԙ��3��6��R@j�\M�����$���ǫ�.�M�*����`�*���3�Z~��8�"�Û���L#��I�&�L�c��+C>"��&>����`��4�!��0����Q菊4�w=��3�8��B
x`��N��v�m��,;r/��p��$ȏ��f�`M�E��i��i���m=�j���a�cϓ��/o���\�'C'j�)0q6�����2+!w<]�a���	�
BG��m��|҄R�Q�'���W��G�=��7��'�۬��H/���0y(�6�C���p�ce�-jO h9᤿w��c�_Q�C��B����n�z[*.��|���!I]����F������m\��Ƀ���lX��x.�-��d�L�_�ϓ �X�<�[������D�p�g���tS�H��8��$���<���`���C��t�ɾ1� h�3h� �8��8}Ր'j��(~i#�`�U�DA ��o� �(�p9�/��@�l���j}ezȋ'�	Rw�(.08J��Ta��٬��e����+�GT�?^e���$b��>�v�؟��u4�]�ưk��=N�jW
в�;�bA��"Z*0AZ\�B�ښYf��V5�����3��
��_6�r�vu^��t_,6AE0=� �����6�!�$�p�T[߾y�H1�M�H��u�j�F��������$���������{�iݣ��؊��;��͡������"i������Er.Q�qŇ��[��$?��H�ܜXrT��*�8�M0 D�{*��ӻ=�NU����D���-��c�mEH�O8C7(�[�7�	�aY_�W�f����;�U�YTF���� �Y	�šߕ��u}��
kp��ܴ��c�~���S~��!�5��@�1�Jl#!Pҡ�c�}(;��POɥ�+�H1-K<J����Z��J�|ٳWg���c�+O%��ׄ��"��?��Uaf���T5�������3P�s�Za����Q`�����)i�'�qNݒSK��WJ ���o4�����u���@ע!;�q`gHx�&?�'��������~cz$q+e'���}בel�,�� Iu��k����3ƹ+k/b�?uS�;@��=���p���CC�Ֆ?���R�R\�����ǯ���8t�T�����d���æ�>f=�|��������,<�& ���ͩތḀд�m���E��&�&�6�2BX��7���[�D�I�
�U��/�e��F.t�~�J8��)�V_`~��5�mi�W�������Ӓ�,w��~�����*hi���cU̶�b"�����ذ����jJ,}�צXR�4l����r�s9{�sUO��+��T����6�;����s���uT�UN�GH!��c�ƛ�@hP���oS��Xx��Σ�&�)��[p�aiӦ���۝wt�>%�P�o3�����Jy�l�(�7ٓ����~�|���.!�a�/�MkI�ܻ�jЂ��oy/}��E���j#_A��@�K���KO�Ӊ���u�V�E�坐�ˌ�����K�P�G�E���r��`���L�$��<�s'�,ӗͣ�.ݛQ�F\�e>��U�[�F3q�������U,{���g�L�Z�+w�L��Z�;T������c�z�
��r7
�ʟ���J���f�:l�IT�78S)�Y��($���hv��� 2�|f����-q}&��&�K�Yb/p9�H렄ʨ>28��Ds��.?�^bag�-��b�.�Q�rK_s^���{���h ��O��zq{�.����!6�{���2��)sb�Ѝ���'�It�������]�B6����B�K��"s\�@r���o�l�)`��Et��o�gQɀݷ�Y�_�[�fQ��%�h���#����!�8)�!�V�U#xUw�S#D�LlA���'{�7}���[ �7	������-A=��3�[����f� .+��J�6�OL��'mm�"��c?_��c���O�'��S3�}��!��ξ�)�=��˙�<߁e*�[o���)@���KcG�w����8��/����LN�K�P�Rf�kTe��o+�E2C�fA�d_"����焘�{�<o+�韙��3�t�QE�u�l+ŀ����?�Q׭����`LĹ:O]��:�г��*U�5G�Ϊ�s-C$�`�=&$G6hhj���M�R���#��M)��x�#RРu�F_��3��D�J�+`�Y�:'3!f��D@��*�@=I�ZA�#�}cL���}K%�$u�r��c��".ž���vb���x��&����?��v���&�%��zFCZQ48���EF�[=T|C�%q�����¦l*�?��J?��� ��iM}��^	
5�k>���IˊV����\�Ajrt���� �P��ta�6Q��,'S#�~ҭuw��>�v3�X�1;*.��=y�@;�`8߳75)�=S,)�Vr}�(�R'r���t^����-�Her}-A�E���\3�@�:����<��5�;��Qq~޿�햂w���?f������2�
U�_D��M�a�Q���¥+�F�A���$S�PVF�$�꣦I�.�hĦB��B,˹E$�gʶ�.,�<����	S@��#��_D=���w�E�@��3���Fu���p�Sn-�+�ǂ��
N/�܏o��Ȝ=�	��l1��K>֥�<ja�?O�O|�ઍ�R��&�P���e1����V~,]w�\<���� �[OP�|��d4��۬�k%XB49�_Ȩ+��Ϫ����L�ZeoP���B9�h�8[�A?�>�xU%i��w�UJ��ekѴ�6�aDS^�
��G�)�Ŧ���<�k˶Sk������R��NG���3f��xU�5e��ٔ=�e�Է�o�A�讻Sf��o���X�j}˅�#��^��#�Y=jRk�0DY�{�(��4���y�۬>^�kw�����#M���2�ѵ�us0M��ݐ��O�Y��LM�V`&�CtYIa*6y-+�m�r�l
N���1����g9�zg�����&�G2�i��PI��B��I�ja���^�\q��,8���e���-�9��x]��)[z�C�>At�����x��Ǧ��ْx�=�*�� B1e\�N�Ѓ�?8�L�0IǷpk`���	��C���f�Y���*1+{w��%��Hٶ��P1�����vS����.k�ER^1�����/�qz�&'D����b�c��^�?/?+>g������f	�:U_�Ǚ�K�4�_=��`���M��t ��bQ�A��@��t;�j���uOu�u���ִ�=g�r����)�P��x�F�:�H�
�Md�
��ܒ�����M/�x<��q�p�#�B_��/�C���*8
p�~���$�8J5��Org���a��\�-��e��Z��+���D�b��Q�~���	���������Secc�3g���`��	�	0��?]}�����6�B�@�85Μ����ͼVPX���K��e�-W� ���S3��*�ˡ��湖��v�ޜ�v�X�N���+���][*O�^�U�J�y�cٴm���%�G;��=�ݎ�!3�(��kY�as�����������5��Ҋ�h�~���ǣ2�M�`�n��)Y޾�tI,��c���֚K�|���m���$@8N\��ɡ7����ZQ�6��OT���_�	б��y����xBa���.�Ct�H�L6<5ؘf�1�p��4��b�/Mc���,>�ut̖;d ?1^���,^�X��Ը��^g,�j=IF@e��@+L'*�[/+�#�I���o��6,�c�E��N��+:.W2Q�@����:��֎�u�W��k+#��D�?K����
Ql�&���Ө��-�ЃA����T��9�i�@��9�;ZZ� Ƨ@��&cY�_%���w:�� x5�Idf��=���'fY~A#b���m=])��H�r�����h�*�x�Z��|"W@��*4m�����n��E'ޏ8fo��
�w�z�;�be��z��XjF�kIW+7a:���,CϺ��5��JU��k�R�B���EmAԗd4r�K��Q$��j�����L�d"+�;;�6�j��Qi�6K��@��-#�t٤kk9,�k��M{0q9KV�
Z�&5ðc+�P��B2V�o)O��k�]�nүk�i+ x&�P^��'R�'3�.�zț��h� �c�؜jW޲��;*p7a�Bz	r/м���dZ7	��_t��w0n�wk��ŷs��G}U�)�cw6�����2�a"W��*@�*�y�NЩ�ǫE�ȟ��Dd��˛W�p�q�n��oP�`tg�U�r����7nбXnF!R�D�MѾ���]Ɉ/���I�-]�b����d$ }k����Is64CK/tO�������)�!.�4��L0�e*D7��Y�`0�?�6LN+�����
�����pYk.��]�S�Y�!�F��w�O�~�	w{fǚ^FoLu:hh>蛳�oO��s��haP����t����^Ei�z��$})�2����
�'�J��P��0Pn����DX�{�'�/�Q�W�fWC ��$z���v7�r94ޯ�F*��t�̽	43�g#<"w�A����)O�<m����zM�# |F����iHh�,ז�OaI�̩7�L<7ѣ8�#���U���,��:�(�,�z6�PG���<w�.�o���/�_��q]Y�g^�����I��/���K�Y����N��xj8�L�?
�~�1�Ǫoo�^�"@h�� �����֘����0��j�{��� �@+O�P�!=hnE��FVѪV�٫�A���}�x�-�6w�L,G�r+��a�9d��Ł��S��W�6�5ȴ���	��1�F�<]q:�7�������)��\�o�V�5�LH0��{g����įΎ�k1o:�r8иwY$06�h#����jwҥS2QA������7���cy��Ac��~���{����t��D�3�"	�w�p���n�fl��f��L*K��.�
>BF`����3ԧ��btV/9?��U{:�^���G%�8�����䮆�3T4�,ҳA� ��h��қ m�:K#p*kًp�S���Q�,k��Kyd�k\����}Q+����qg��a�㦭:��R�⏣gV���`�f�U ���+ �-�HȔn���/y��KT��C$y�p�JX~{
��p)%�dN.�)�t�=+���_G��M�C�k�r�9�Um-V�	O��%��~xdh��;֪c��ޑU��z������^���>c����(�T}"gvG��3|sƐ<�c�G�ɚ�"q��)3�t������9�h�?�g45�M�H�@qEe�_4ZMŊb���fF��"eX����>�8�4���y�嗕0���~��)��
fKⴥ�"�������#f��TG��tI����P��Q^�WG�F��:$P�M�kSAg1Z�2�q5�ǅS�kX�yH�U��^�
内E1�F�Њ{�����7�?
t  ���):�J�t/�˩���A�y �䠅鍹��[��.��H�u��f�ѢSw3-���-�,:1��+�ǵ�Ť��B���d�,^�orh�俷F
e���E�-:�����ry����V$�B!�'��*�%B�\�ѩ��m=Of�E? L#N+�T�v�=���;M�c����N���H�$�t��)�*�j���.�ѩh�8?;�~��L͉7�F)F��S@���w��;�H�v�],�Ώ�D�6�y� 6k���C�=fԒK. p���}%&��4�J���V%ݜ0�,�QóB҃��"��pԉ�o�������Ƭ��!m�	�S���L��+��ߝ����"��,�N�뱵��"<9x8 �F�X�9#�й\��pQ�J�+�{g��mP�G�����I�Ĺ�x�F�6��
U��M���?}$�1�`�j��<o"�=��?�=�e��C_���|��W'���^�FS)M�ņ�%�����<:�v�"r��rue�R��D�����Dp��p���AK!�(B��(��n��J��E�|.bP���7�0��@���xڲ��iL�ݍo�ڣ��1��Ɋ�{�Ǆ�v�FXh:ڜ�F�n��Gp��I�;���O?�\�V���'�yQZ�J�c��S����>wâ-v׉�36��ᚰ,��_�1G��?���F�[��D���wG0ф���*$�]ў���=~���j�Lp�6A���8�7#�-�r�~�3��v�s ȟB��Kn=��aB����]̜+��D�����Bs�uk���c�_u�,�����ƞ�gq	2|�����y&F�Gt���5y#������׍+��Z&���W�6�}��SvE���Iv�5W�3)ȱ>D#��,�g���� :��]���ՙ�������5Zš�vK��
����a�%(b)���Or��?{����z
)�u��� �e���ج��$��c��o{�gð�[�\m����i�+<x�c3��BdK���
����_^���t�j��2��������l�$k����q+�3-�"k3��N[��(���fd?��C K�<Ԅ��A�=c�S}{t3~U&<�T�V���o��%6�zE;�#T�a�����l�[Ƣ@N�R�ؔ囪�~�4rn޷�h�������A���C~��B����yom�NٳD�WX��TN��C��j�.\��^E��8��^'/�q.��A_��,A�+r.�<�@�Ik5���1v�X(E����>��>�[�k�Ҭ" 7q ��@l�B%r�yPp�2�{�A_�
�I��;�7=��= �QlC
_B;G�4���ȼ�Sf���)�G�������t���*8� ���}~%�Z'�Fm�b���v�>�7���`����[�v�aS�[J�2T��x�CyK����P%�� ���l��zq)����g���7�=jw'%�R���O�'�=���hM�\[�r�9k�?�a޳.�m�+�6I�(�J��n���(z��>
=ө�z ͟�;7�ȍB�b!�;毂�����tmj�Kȕ4��p���C89�B�H�C��a&� X�&O���֢���u�rf�G8�VI�V�B�L��\�=G=k��ó�	�/o	���(�I��9M��ߏ/��r��M:�hխ�c�'86h�f���"J+	�0O`T�������+k�uTQ��a^p�Y�3c�� O�a>O �7n+�O�����ùW˵�\��W�&��\�!eޞ@��߇��k�P��͚ܓŌ��>�{	�j�D&�s�Ѷŀ���x:�9*'Y%xN��]_̝-�~b��%���b]W�ծkd7��8�:|P���8�<�Т�콫9E�)0S��&g�ꊬF�;��K���bJTx���.O�|ep��$~?NU����gژ@�E���~��Rd71��|�?1�2��'��V��?�f �0j9N+wR�4�*:��́t�n8ng��jo�(�N��s*�xG��`eUʀ�,���9����3�9{P�Pc�x7��*&;w�̑2�tNfk��?<(!�dӺ|�t��A=��"w���S����������fP�YG��+���Q�N����;$�vI�%���l���D���m�6�O7��T�HW:��R�g��ْ7:m�� J��oZ��t����F��;��vk)kߜAP0�1
� ���r2���=�rt\�a ��z�W��h�SAYV	�����\;�Լe�:��u矁�Ѻ�q��Y�$�[��M�k8�����2D��=�i������ k��}��A�@C���k-HVX>��h�5�{��6}�ڇ�N7��\���opUږ���k�f�-��U�:����C��;��\��z����:Q��-����yef�ƶ�q�aMma����{O1X��$'Y.�^�R����<���(�!�2�{_�T��9�rX>V����n���K��������I2o�:`����Z��确yHݫΠ]C��<B�j ��B��al�v�]*�7���_46d��vq���C�?Tu��c��Ze���RD딙��8��<��GzZ�y��W�=:��5~���f��G���5�cK'���K���!�I�6V�=J�ӊ6n[��#9�����Ϡ[�R���k}B�3����i4�QԂ�P�����4Zؑ�-%��ʨ$��� G���)b{��>��9�/S�c#���S�C^�pmYv���?&������%
&XH�D�/}�~�f����:���-�����)"!�R��g�`���gfg�ٸ���L���!��ź� ����F&[��Ӏ3c��f2��+s҂����Ϙ�b����Ԯg�_1�uG�~���Ʃ�qMw�Z�3x��������53!�4���R����Pi�o:�)Q�턂�4:-�U~:Qځ~1�`p���[��!���Ƴ�| �W��dR4Ñ��o���Vs�I�z7��E�h��A�D�� N�}��Y�o�2�q�1+g��0��GE���&s��H1�*�c��`Ճ�p��W��%�X��6�����E�y����r5=|ԛ
�w�Ij
gR;��#��B��>=z�tq��-�U7^m�#,x;��D�Xί��@��&~{s�$�*�EG�bf,���;�!���c�F��A�KG�_�<�v:b׏��ō7���r����*���d	��+e,��O�ɻ0v*��Ȩbol��G�:����}�}������#��� t�jb��4ާ�,W����SL�p�c�c��bM*�K��M.�qp]���K��sO�h��UQ��8�V[�tr!�O�>�71dʝqk���v���G<�ݲ�w��G
��!^��T���M-��7�����_�P6��A"s�N=!��5�0X�l�R�e�+��L(ץK;>Q%%���r&a�<���QUsL�21d � �	�j@��Hd1�DG�V��|,a���QK�C꼿�~dM��o�ȓ����١#���;Ca���4x�wH�B3l�,s���H�v�{U>>�ڶ����QOҷ�dC��P{�]40��������,(RM��mn8��~�UCrb��5a0@���g8�N��&૪d��{AUP�^b����CQe��%H������ l���7j������ݘk>�����1K=5���4b����/ܮ�ԡ�A-��r�����:�&qw��-1��v$���O�8�w�l�O1L̓���>�T<�$ +lU�X�La��.4t�F�]m�_`,t�L{D2^9�x� "�����T�!\�A� >��B^w��^�d��</�:l��10L�z� B�4��(��8B}u��J%�[R��}�I�5�lʴO?��^���DQ��&L
f@�aC!H�*,�a��F�����kW�w	�+�נۘ�BHa�AAw�� �~$�� Ei<;�-�uM�ӳ-��>��~�t+�M$�F�a��T�S��F�p�tW)���BPb)6rbC�Zy���"�ǡ���u���6Ag%i��n�	���z�6�US[�3{��c-�IX�
�l���]����,��49^��O����V�l4Z����D��0d*A9�/�=!�&3�D�K\�
�˃�oNx���+��7��;J�"��S��K%�\x9�
&��X�z�1G��L�ڶ�6�e��5�9i���T���f�zp���|4d3s"C]w�'fK���3Ŀ�^7_�T�A?�(�ZY��p�?]�ij���k?�*Q������G����]r���Q=�����5���-��.�6��S{u�Ob�UBZ��+�u)�Bl��d=��l���Cu/6A��ۺޟ��Uz�{Ń�\0�<=���3�I���z1EH��{�+�&��USiG�O�W�=�uY/�>��ߦ�JM�M��)fK~��\��\��M�"���+����ο6��fb���pVm�6k���G~ޯ\xS�)!)�k�Kr�-�+�-�ő-1�(���"6^�̎?�'�oe.l���#��.-�-ĕpf�}��^Ġu�6�"�Z>q��2n=�-�R�pH��p�":Cc���U�Oo����V���
���8�n�q��y^�U=��8�$P�/f���y����<�3�u�]r���۞CO���
S��o]�p�!�Hg���Rqo=�ݲ�=�����md�p��g6�c��|j���պF��tW��Xd�!CL�^��&K��D�m�o���%���A���J~OA"z�� �]5؂���8�Y���A�P��t>`G���m�Zh����i�t�b�Y��c�S��i  qؼ ����	��'(x��EdN�޶�eƩm�2e6nr�ڳH�y]���5������g-e���-�韸��:��m���ҍKзaw8cي!9�%a;eE.m�M�����{6Տ1�l��y���&s�k ]�I�"�f6?E^߸��ɚ���m+ݪ�t/vʀ!��a2I'H��_��{�*���L&�l�*����p�+��Q�p+e�Vh0m�Χ�s�Zދ#��O�Q�mSN�?�VF?)�!�J��{����Q���\oT�K�j��KY�ɉrܿ��{�+Y�ê�~V��zC��Eiy5�=H]��
�7��ȷ�I�66V���y�s��]��o��܃�n���c��YN"��1Iv��":8��`��Jy��5t.B���B��*7��.hJCRĥ�&���]��<�àc�M
f���5b��d�mj&m���R�Aߗ.�B�,c����El��u������dљ�ݥ���"%�!`A!4E�YPk�v>�\��imfhB!��\�u�Kh�I%��Ip����^�a	��#��l�<���Ӫ6r:�5�����8�N������+Q'M��o����7^����$����S݌�X	��ݝ�����&$$%�U�h>�q�%kVU]XN"	�z�{�v�F�tF�Q�mr������ ��V��y���Bޅs�8
�3)���:����r쯫^'�%�A/�cm��|�q;k�&}E�m��kw��F+��_�WKﳙ%��5-��.ِ��s���o�o�P?����pB�U���/�a\(s�4�Z^���/�Ex����+��r^��=�l�L�$�qȤH6��9m�Ms��!�ʳ�!=ս�_Uˊ�<7[*� S�+�e���k�G1�%�|��>�����<SP'r�����#b`�����v��)g�V���Yeg�z���D�=��s:��r��^��D�2�t�,�Ӂ�_���b��{�z���'m���ןJ�eu�����a�gۨ�\�EJ���d
��^Za�� ��8|n�ŗ�a/@U��H�9�|x@R$�RPu�jyX�	���13��3[&("���zد��\�6E��`�)C��݀E���5��ڿ���6�d���I�A��XB��8�$�W���e��hc�BY�2�Cuoy�a4bFyHdH�m��q:�����A,�����4�������׃%�H膯��)l�~U�	�}NP���~L�o+�}��$�c���;g�5Q\�ZiI*�ܩZh��c��i�$�ǧ��AUj~j]ඎ7�|_��u�f��ֺ����=�j ~Ф��ezj�(x���0���:�2����&ճ)�ZC�ѐ҉�!��G"���<�f�r�1y�z�8��ay�R�Е���|�x_\)��]�d�WlS{?{T77�^��ӿ##P�oz#�ҝpCBA|"bňϲ�4J��П���UM�_ן=\J�$.3u8����Y$,"Z@/����|j��m�-����KKOO�M���}5���7��Nb$)�{r��冀�� r���w�9(iF�i6�0���y�Z�zW��1&�Co�S��ue}� ���V+��5$���(I>��5NΗ,n2OLs
#���e��x�����C�X����r<���Gs���4÷,2~+�+iH9�h��1 ���S4���g6 ��n��1+:�g/"�J?�_co���:���J_2�1���A�U����v��EXC��مۭɉ�I�Ո,E��+���}�҆]�Q`�$�*0=�����s�]����7�����l���5 U�����rz��g�X��>A7Q�*����\ۑ�����߃Щ����.O������vy'F��{�6q=��+����e{���jgV��У���S�j�q��L�ZQX����8E~3�p�	�(� ެY��_(�c�B1�;dE�.t���l�i�{��m�>�z"��d�F���l�X���ֈ��M��嫍���2YjX=P�*���][�R�K�0g�r�X��p��y�D�Kt�W}�R�WQJO�#.��ڄ�$�0dw'�-�`\��dpk<����l�E�~��e��E�<���N7�%[T$���K�]��]<�7��/	-RM�
bZA0�PX��E�;o�@�v�cӫ��%]`�u.0�dO�;\�@jr[(�t��ċ����q%�Sw�2[Zw�Q�!0(�[�Z��-���[-�3�\�1i��e$��G��u32.g���Sw��,�wA���5�^�H $���"��!������9Y�z?'ɧ�؛_poT�2�����xII˱��������ZեK��L��-�1Y���/l�;��c�/�ʘm]���W�%�ꧫ����6�5�h,�`�=�$a�Á�:�$�{N��7k��Z�Yٛ�a�D<���e�r�E%
�/��Mudc�������-T6<pF��
7�e�#`a�䀕����v���]������XP����7/�C���k�:�Р���(���C������,��0
�A�����uv�U5m��K��~d_�3`�*����߅�;4���0�)i9�oty	p1!:	.�44)��.��j���U�.�BU�N'l��͞�?���|xMP2b���{�*��o��i�������<8
v�L�&�YĲҳ���,	��A�E
0�b��J�5t���M@��,������u ��̣�����}��"u����*��u!�'���Ω~�����WQ�<�>��B���/�ci�~F�p���k�s�'�9�')䌕stǹ(Y8��i��Nh�ã����`㣜���E3�ْ��_�8o�_��Z�b} ��e<����\,
)�pi:���KU!���"�0�/��K����Mp�m]��.@K��V�~�E��j��'�Ji�y^�g��Z�F��[��F�!�hc^�K[�����	�r�ob�����9�M<�,�H�̆Qx�Xc�����pǙW���ⵃ���n��
?K�=���n��*��p����;"+�t>��|~��՝	}to�
�rKT��-x����?� ������Unw���e�&�����la�����_ Uh8��� ��f�h����}�rpH/s�]U�� x��I�D��DA�$>�6vE7���̋�	"����Hw�@J	�%j��x!�>ؘ3p(nqDV�>^4�7������'��L�1o쉈�ƣ@�Y�XF���@��W&j�����;�F �ݬ/o١� =�6Y:^k;"^.eßd�^bՌ��l�b2cǄ w�a ���1�Ղ��DP�I4�`��H�Hpwnş�O�/�w�i��j��Ϩ׈�`X�%��x�6\9����F�'��Ǽ���m�E�&0��#K�\v|տڰOz���o��xu75.�Oi/�����[E�dL�!�өW���3�&��Y��f!�!��,^��^U${��t����f��hH@N��V`� ����%�0	��q�Y�k�}��/���8�N��s�<�fz� [�n8���� �Z����V�'�O~��tp�m�3�k�����؊�1�[GTsNu���+�KuI�1|]�WZ��vK��)��֍a]�����U4�F�[��8�	��z�K�{�|�a��	 �D��/����p]F	����8R~�c=!�e�+	�e�j���֨X�tt/����5n�u��|U��AbGbY=k�����Kd��mY�4o��ŭ�T�"C.����Ag�����Puz����"�j��h�vmt�rB��wä����D��Ow@S���)T([:G�$	G{�	�r��V'T!��h�5L��oncaٰګ�/���H$�yLl ��;LOq�7^��7vݖ�.�|qe��������$�6���x冱M����]�RS��z�!,�+�C���7Ri�n()�D�@1��>������Н,e�������K
��q�<�� ��c,g�r�N�Z���!��V,�+����<GQK���9GP|U��ԿlD�D���	��.]�:,�WP����/p�b>��3̴N�m��������3u�/�nU�5bq��%cl�O,z�B���)�p�H��fps�{���-U��� �I%0�sՇ_S�yUO�>��"/�?Έg3�&��b6l����}j�������־$!�m�!HZ�ap�e���������D"���M}W9��&btN�fS	`�;%�U��yy+��/���&�4`Rq�2���?V'R� 	�)���4Ly[�M�h���eMG����6:)�C�Ⱦ�`p�3���s�l+�ϔhq�+�P�FaG���W!8�<
Q��Z�H��/���z(��1�����y:�@��@�4sn�˲�Ck_��&\}[��^j��qM�T®����bޣ�2��D3S�,�T^�l2�H9Y�yf����ȍQ(�O�~	�6�}r��jê���̼�pf>�l��~�JB1q��#�Q�<�1Yd�ٛ��|�Z��M���
'\$���Rv��`�&�5���{YW3����7��~�Ao�{q21��������@iE�V2K�uQt���,�����g�Px���v��в��=E����~�48�W"(�=����!g���t��+�nbTӾ��X������m�=��$��N���z�ԙ_��~��#���y;5%e�B��#55xsM�Ɂ���I~T/���Q0�ݧ&��i�˟���Ԝ|�U���ܿ�[*�Y �"�G�3~��CJ��Dh�#]�ek�m�Ȇ$�n��������R�&��AL��XHd?��سq��dMc4�ɚ�Q�dʣ�~i^̠�SZ�S�ƨ=���sȘǪ�)�J[cɺ��[M�I��N"֙r���[�d���߂9R�C���� ��d1C�ډ˷�k9DVf�C'�u������`���3��賎�	��җ�f �|�)����9ǵ� ��+��Rl�F ,���=?Eb^>��n�[��x�L�mS,& qaPP���ƪF�z>�fay�����z���<n=�E��	��앜��S(�g��8��:d	��P�ڒ�v4WZs���Ŋ���}؃���U�%�ӯ1]����������P���B_��Bf�0!,]M#Z���!c*X�mq��9�_�����ߪ���;�xbh�L�= L���f��Z�����%CE;��ԟK"����������*r7->�Xe�Q���
��k�V�!�X�Zg��K�����d��Sz�	���굲N���Xv�`(o1��?����~-@A:e��)��2[�F��u�cO_fq��ӕv�0�L/�������O�S4�ҍ�\��u���"�o���ݗvEŷ����ǏM�Κ���sJ���"�m�70���(�'� �R���@@��6�0�[yt��~n07�f��*@�͙��F.�yޖ�c2�!��o�7���l"KR�p�(�fMԽ���< ���I#}D��߮�x��^E�M`���M�ݮ-a/��G5�%YL��\mdwt��Sz鬛1��h(Ud����� �/({�`�|�X�a�&+������mOV,"P�ǿ�Fh�Z�Ko�X?N�����H�A$]\����M��e"���+�Э�!��S�7d_�oW�?�����x��<,4�~^�et��~<~$C	�][��{��<��^���_�/�?K��mm���S�>��rI�)���8ċ�R�Rv<������h�����hQ��t^�#d�tK�hSe�JIu�>� �j�bIta�1k�� �o�&)�������%o�L�~n}��9=1�� ^(�Q���fI�Jq2AT�A3G�y����V
�N�xY��QWPx;m�a��*u��p�5�f�#
QyM�vсh	}��4h�q���L��J��:���$qE��1��p�i�Xm7j��w�pԐ�>9_�� D;�eY�ۇh����+�G�w��!��4��z���4v�j�ڬ���n���m
D����~��Co�b� h�!��ު\�jP��W����ETb�K69t�|؁;0q���̟k)j7#�R,��'��]_&�eK��9Jp���z�����Y���}��@]4�Cv���Q��B��Ցg��h�*�p���n���N�9�d����S�/�-���.��}�Ǘ�u!���D��˝ϱǊx�7d b���ı@>#V�����[�྽ݛ���p_:����������1jO��F���ЪS�3!weJkZl�WG���U���\���Q�c����Y��ła�i�&k���P.Po�8��F�Q%P�L��7)d��p�R|�,��v�`�V%����cT�n��_*��p��͵�]ZP��ȋ�!R�polX#��H_��>�L�{{��#���N̺�ޚk�y��� s&�Z�H�|>A�Vn2�KF�g�иRZ��A�?'�4Ȫ��J���bFy�z_7��ǡ���:]oڣ�(_�iݴyI��!ӈ�㲒�>�[�1*�6��[Oe��٧��uG��y�xI�mId���`N�Q�A���FU�b��~�|�u�_$ݏS��ǤI~��z䗣�p:k��������%�g��H�B�H��=t��)�x���H2�D�O�4Y6������PҐ�"x4't>`�מe��ɲ<!u��0�:�����9��G�p�~Z.�;m�J�k�YF��3R��c3�/��t�s�	΃����ݗuZ�&����1����;��<@x-�N�멓�����t8vM��/{�UQ��P؄�� �WE~tU����̫�=���<���[ka�qn�h-w����q�#
�P��]���&���L��٨f�������� ���߿�����M9^Mgu�%�#sD"�X�w]k�Ѱ�Y�>����o��۔C!1��x�#�4�3�4�zc������L�j�X��� fn��0NE�T'� �&��RMO���y{�z�Ƕ����6M�J#���*�lj��e[���ĬI�B_ޕ�}�P0+�aao)�95�Q�!Ռ=����Q/�C�v���۝eӫ�֫���j�\�6>L`ʼ��1��*�t|�4�st��SO4�B����"���7��p;m�M��8�:�I��b�t�&3������ ��h��+��-�(���G�(��i�^�!
�_�4r�t�{K_��	->��#��k���J��B��^���v�#'�ơ��q"�������]I0�]�:�Ր�w��&"�x�?�0������g ���@�z�w�+���Cq9���`��9�v�_�+G�܆�ۧ^GXK%r-kЪ���������(�fڥS�
,�)�oPf���6�Ek��څ1�;�:H'+ea�D81�lռ��I���;�qӚ�^N����e�,^G3�_��;�Q�&@���&���X/�j���Y0���h��c8�yF�Ӭ��"YM2�6,t"S�I$��r.��<`(��s%��V�8������=�\�ON��B�1h����GI%�������O�2[�V�����Gv��[�ٵag%�;�``�h>eu��Ե�[���n���Ƒ��ڗ�K�U	=���]w7�������/�H
ßz�u#��/����#ӻ�tt��?r{N͞Z�8dk2�ڇ�[Ç�~�6Hy]��$e�ZJ�9oBH���b_R�Q8�x7`�p��]�iV�T~�X�L��GЭc�!g�U����)�@���3����Cs� V�+�oF��J!l"�<<I�,߰��m���N}���K�>%ΝBS?�A+��t��6u��[��vM���i� �Řpq�4?��� ����$�{a�_GO����d��@?�J ����4&���L%��Ŝ-W�=�����_\-F�5��}�%���F�w@Ը{�W�b�P`�>�~h�r*X�Q{]���+�Ђ/}@o�V@�"t aNd3 �/���%�^G����+�;�]������܎r�/�������_&rs����F���q��s� �����f�?FA��{�����@�tN? 1t|�H����/w�=�<��}2C�~�<�1��6�v݉���`�W����?4~O����~��Qz7Sş��BZ�|��F$�<��87���w�YO҇��8�a|^�@	"O��+f;�>�<�ǩ"���k!x����?����&�/뷫1�}�h��˜�V��+����Q�"Z.�h�,�%O`���������8x��^6��o
��������������Rn��%���p{D,�D�T�V{4���d[�&�/�3l���T�M�D�� �i��m��*�Ά}��Q��)���4�^t@�����ԑP\�}�i��-�h'M�'$L/���@�ᇑm�_l�a��`�SR����5|U R)�_�F���z./j3�H���p�"��~���K{iY�7���@�yc�7�1W�*� D�Q�5cC�{���ss^��5%�kbT�rU�Tҋ�q��f�!�)7�_��"|9��"�93�Ǚo��3
�4�7�O慀��(׭&W(��Im�b�;�?�O&}�G����Q��˕0a_ǨxY���BI�� (-&3	�nv0	�`�Q����m�qNop5�ZK�]� �7pFx�L�M󤽃�eb�`a�N
��䖊�M�R V�M�È�}�~D�m �d�l�Wǘ�N)���$a'L!5��ڞ��e�hhfP5�iZ�b�B����ξ�)����e�k��5�7?+�8��w��Q�#��w[�m���L�?a�2#z��V����}��pi�6���)��SK�g�iT\l͑nE�]L�PT��!9��E8{u��	ο�@o94R�߈�Z�הv*'��Wlw��A��0��8�k�W7*�?�Ă��1sŸ����<�9�"��V��$���UE�Ȯ�nP��_�]bZ8� �'_�)(Lݔ=�¥����ʉ��=�I��u�j�1���z�sYj��Yl�0��-��*�_��f��,�ӎfT�[�����n7���{i�f)8�.��|x\i
�a^oe-�X^�R%����<�YY�1�G�=�CV�볶���=�����M�%���D��rǰ�����
?kJ�f,���]�_�#I!���P�"��5P/�R�k6>���̛߫�2ߎG_�4t�g�ϡWs�&��~��8���4s0� �%ۻ\�\���=� #r�&����h?]��&]���pP���+�=[U�����7��:ߩi9�0�m���� �v�sw��oc�@��ͬ�"N����X��G� '_fS���$>4�~���S�t{%��
	�z��š��{�P��7�f���􉳱�QLO�}���(�"װ�N�C��Qx���[�&~Sm]��logY�Σ�a��}��P[�]�JR�G)�r:��e�-ˈ�F��}���Њ/�j2���\��:�_�}
d3�ܒ��o
�(�rX�:��H�ϣ�@�98����W�����������iIO�p%%C�ny�If@aF�"fD7yq.��E�~��`�b�h6[2E�l�Q�m�^����ԌSz��R�H���.<Õ�7�굿��ˬ(ZD�Gt�x����*<��N���d��3�G���g��(�H�8SU0�M�l�[��%9��M��I�(������$�kH��R�{�2U� �ҫ�]��+�S;/��ɴ��/�0C�u�9����
�n�P�m��ReWtNc��J�<����ި��+��jqڤ�2c�3#Ty3E��T�y�[�$�(���sҔ$9⨍�ɠ��Rsپ�Z��+?.+���2�Ѡ��� �4�_4Rk[r	�ݐ��@u����L�z@]���+p~{֨ja��I��%�qb"�'seD���]J���	;a4W���Z9���}�bUe�Ll\o��Y~'�y�AA�\؎����d*TGG)����D�C�ތڑ-E(D�#��w�!63S�p�m�3�T7�;����O'�Y���Lޔ�~m�d�RC�~Q�m�p�O�,��Tw�갅jUȷ|1���X�iJ�7���F\�ұ�G}��z�v+}Ȭ5@`&X\)>a��w$����&�#�Øъ����%��0�p��6��å	6��#��+R��}�
oIWy�Z��N�ǈ2���ǿ��'~��&rA�����|ǐ�;\$��BQ�y^�`̇0t0�G��m�H̀��#\�Ě�>�>~� �J?��<�`^��5�<muU�:T8jufu��%s_vK���?
��%`>^�|+`��<pjk���/ 
z03F���V=ΕXl��3=�耉xq���e�e?�I8�(ӰZ�����n]58z����ټg���$k�h}�k����䠸����c_y����Tw���}Qr.�[[�p�����|�2�c���VQF��-ȱ��Η����'��Q���_sǲհx�44ȝ,!�`V���W)Wj��{�E@®qn�Ʌ�[���eb!'NՒߤ������o��c_�j�y�i&#֯�`�ӟ�T�����tU��R��N��E{� �4���;���N'	�����V0�y����sHvS�}mAx������G`}WcH��ɑ��|����AIR{����-Pj��I҄�ފ�� �z7xU�y������N��������%���,&�{4�SH�f/�2^��q�7��Opt�(�6��\"bs1O8�� �$Q�ȋW��yŋN��k ��\�x*��=��c�僳����˛}��L����R�O��.0�g[8�ӑ"_R�����.c�]<H	��w��**,)����Rj��9�s��rh�4��gK;��� '���J?�,�0g`�kgo�w�1�L��� Ѽ����t{�٥*��`,��[�Ur�'��!�R��m��s����h��Y�� �dU�G簃��5�B����e��<B���]�J#ڀ'���!���ʽ��q�q�"�4�fs?��7C@>c�����<F��n�.�ޏ�_�_1+^'��1�à���9�ZO��M��q���Ӆ��'v��]�J��?<�7@�M��P�b��Ӕ�Cñ.��SXa��6V`�4��5�$�GL�μ|�qx�E����U�|��F��ہ�*?���������ܺ^7�.Z4��e�ŦY�@��G�|M��6�~�ބr!�P�PF*�1��Qλ�ٞ�}x�ʏ����u�i����_�6[ ߽ͨ`�t��_��a���#��r�h*��^�V�yxh���gDb��3��K<���Ha�H����k����M
��˷�A�<�m���&��6..�Ș�Oj3{�KvW�1� ��C�<gh}J��c���h�6��k�,)�^�ax�z`�.3��^��ےPY)�e�t�ٮ��WU��c�_�8J�&2I�	�6=����FBdwx\��Z'�����$cL׮j��S�ьZj�bX�\|N2���OsD��h/���~j�9�(�̇�O�����Y?�c`���bm�U`����VZ0mu��s3
�⤰���e�o$GC!jX�P�jH������=�&�1%?�NS��s���ܢ�J;@�P07���9��n0��c�ͮ�����-�ڑ��@>�l�: U"�~������g�:���C��:=q*�IKҥ���J���z��$ƐN$���wA��HK��3Rz��y��ߑ���~��8�;o���Y�� :b�c�ntJA�w��o�n���E.	��Uu�I�gF��b�,ZF�\Q�ѫ��/S��ѿ-z;+��:]>����k՘��c`���e@d��R:",�e�֫�lv��r������}	��x�7b��ѭ��mL=cW1�H1
���_�9�I�u2sP��f��Il/���C�؂�8��rB�O���SzԼAt�e�?)(�N�g(�2+���0H���#��mvu��}��6S�i�a�"߯�%0 ��Ф��7+4��-�V�f�J�f!. 2#�Á��SSX�s����/���8'͏�4�K������.\)IN�a����,m �-��݀%�X�c�+rP�^�ʾW�s�L��過��1���bY����$��/On��*X���l*�H�ƥ�hJ��Ȗa�n����m����[&1�n��d^��n���^�Q�d6e�����K�����"�3W�e�߲K��lZ��@mD5�1Y�\����ӧ�pA�WcK8����	�I��'�}ۻ����4qJ��d���I�#T��������IE/�n�e˶��n+R�p_��ȋ�ɇ���-��#��(��G�&kgc�"&�~��"�������q��)�~�`�9f
f���+:�ʚH�Eo��.~Cp�ك�򥝂�5��������r?y�w�B$���J6��'���\i����S9��Q��`�ܫ�\����F��/ɝ��:Js��}�s;GhGW'��s��?�`�%|.��#�z���k]�3pT�4-�������o}`@?�^Yx�22ea�M������-}Qu��F���e&d�TyP"	^>���%�.a"���oU]9i�q�a����F�%�j�q&`#)5/��{���<��01=#����H�w~�S��,C��N�z �:�t�Kd䨀�t<���Iw�wI5-�_�Ȩ���;Y�k�9�g�@^�E�w��݇�sn�V��^b�;�'%��+��!t,xM(���Xf�v����Ü"�~�X�P?�>O�za����A��a�7��,�:ms�����7��I��*�+6��Hvy�wp�y}��B8,��_�7�(��"b����1�+d�bfL-!F A;�jr��d��֋���� EY����0H��H��L��:��3jLs���hK�7]�ͳW���
�L���OBȞ�M����Զ��k��\cJູfⱍk�/	�����=%�`��dKJm�O�=y����)�TW$���}(�90��U�7���	�g�6Q�������ޖ�Z�c��l�6c��'����F�Ԟ�o��L�����?�x�n�XƜ ��pJ���������$�0�
��E��N��.�����nU��T�X�U�l���~U�d[�E�
x1=:#��|\ �����Z�����e@�)��u��5PO�՘_/zp�e:�+~9?{�/�D����(��tT����%��v�_�U^Ί<��/�d�̢��ʂC�gC7΋���ZU�0�xE�2���S��&�Z�6���w�a����DH��z�@��?�L�C�@x��f���R[�Y�0����<�jj�L}����l��v�\9�$�~@����e#�"����b��A��{o>:(�>/3#G�����9�$)�ڔ��{��,�9	@N�1��'.xaE�`���$*8]y�L���<� EX�Y=�z��q7Y�AI�e(��=B� �P	�B}�F�~/4�����	~jX����c���+��@�L���u�B�/�KYm�KN`��]tf<�[�U���h��\{�y�$??�C1�Iw�%�������V���U TO��?a�O���OC�U�t���8W��c^ۻ�:�@GȪR��`w�q�]�Ǜ1ߴׂb������V�H�ր�#b��	�*���:��Cz��푱���/e���n��o�5�?��t����E�t���к��~��l:W"3���"�C��q��h����}�����{s�ף�	+W�.g{&��K�*X�oEC�����Ŭ�=�b8�Z�=	sJ� ��v�(��ly����� �u����R��.r��?(K��/ɟ�nZ���#�S�Vn�Z������ C��XJ̜+~h!`yY��ӅBY�����%��g�iC�K�f��R��fP~�1=�&_t�r��z�����i�v�V���8���f�_�����J��A� ~�1� � p��uy�W$H��@�&$�#�YZ^k��#����veɵ��#-�|#����	Z������\r�Z�lOO>j&	�y(��4�Q,i���
�������"B9�Ч��9
�7v�$�@��������5d�΢��S�����AM/����gwHJ視��ǈ��*�EZX��+���\��T
B����(G)�,����4e�s��n"��U��w���`�N ��/����ژ
��H�O!�=)óg}���b���M�����V]e�ZT{\��p�i��)��Y+���fW�b!�H��ހܘ���ڂ{���}{+E��������6E�i�3J2�z�&�u�S}@�e��G�RLs^д:��aK�>Nm׫�,C�ͻ��4g��E�z1�3L�rW����?�z�e�#��_�婦S���O�؀��u#�9�?�#j���σ�O��^��?�'��~�\����h��G�f�����G�����9��
]w�2(��,��_8Fd4숱)��,
�(h�Uz�����}� ��ۉ�iP��|��S��&�0ne���x=Έ�ò>`�d�'{kz����p|�׊�#7V�П(�>�W�dԷ��C�~w�)k���X��P���]=�2?����G�$���Κ�� oARY�1�ALyGj�߉a��*/�bd�]��A��!S���8s�	�n�n��j�����d!�F��MT�vQ�Z�nܜPrꓱ�X /!�2��Z0è�$��4��]R<�ђ��d�!cD������P��A� ���f[L� V�E�Zd^�L��%JWb���@
.^��,/.���#4���uPNg[j�����~Ӭ��r{ޑ�8O�8��dvZ����2�X+���IZ
Xl9�<oI4Ԭ��������	z��[QG''ë�Z+��E�,�2opF�C�ٰ�I��lY����q�l��xx���Ǯ�>
�U8��<�0't����?˙�t�X*%�b'c��Ґ�4��L,��x��rs��vҮ����J������M7�޵$�Q�nZ}T�����l� 6^i4�D˟Ҹ���Ȩ� p�>y�Ñ���"�u����C��/;����^ֳ���m�%�p��o��d�~g����n���l?�as��Q���q��gQv�*+p�����a�"u�\R>{�rxM�th#:X.Vъ9]��N3��3��w�v��j<U�5�����6�����Њ2�a�'gd�5��;�0�$�}��2�P��A9 X8I*!�p5*iN��0������&���T���k$c����fg]c��I����U[�^�agȉ�_B'��U`.^���(���:�!8������yd�@g=�7E|o%�����T������8؉����"�?<��cn�QK�A�p��i"�H�Ca�9�`�I���u%YD	�bU���w��b�I ���`f+�f���$����4�8�֓@�թ���65���5��<@6BZ��C���� �&�a�w�z�2������Ӛb8f��D������k�k8޻K�Ҷ�bD�(���O�f�I���c6v�_�k60�/H��fsSN��n燪HU�Pof��Tk-y�@1����򥢯��BS�؀ݣڽ��]�zS�x9�=ǔ��}�1/[���p`?;��n�4��@�K�we���E6`�n�(��GB������&u����KѦ6

�Y�/�
T�7}2��m���E����(H�J��[��#jz���<��n�wm�DZ��&�P��9�W@?N�=(Q�'G�V���Ѻ�I=�ĝ�x��o[y���Yf#��5_�gj����Ď��2$�}-$��}��[ND�wQfv�Wi�=S����K��j�n��,DU���3�[�W0�P��b(r���7�CȌ���*
wJ9R^��@�t�ŻBp��F��g�hI�T��q*�����UY{�(�w��Dt��{���dj>�j�	�	TL�.�b*>�;��VuD=C���� E1��k_�p4W�K�U�9L���"���Ұc-��K�TiP�oh4��Db�+���`<E �ehO�GI���Kz�q�0�����1�.R��N�o�^���Ŵrn:)?0?`���$A���6�r���Ԟ�'6+�N�8}�n�
g��٨Ұ��6�0{tI��Z��)��"��mY&7{��י��!�� Fj�[V��/��7�n���Gh���V��D���u� �$g�u���~�$*�ө���m%��L���{�h�սg�j��vZ��������S=�w���
h �Me�e�|�\W�&UodwUY����q̙!Y�yY�|ŪT�����<����T5���b��[����Pa�&hwؒ�%�e+�Lr56���]X���<5A�s�x�,��+֯�G��=������ŭj��}���R�M�����b��?�x��)�}Q��Kt�L��c�IbQ�8�B��zȣhi�>n���l*��{8|�,����Y�j^@aaT�J�>wȷ���Hb~yLͬ�?k��7��.U�Ǔ�7�"�^5���J=~0Ύ"�}�=�ځ6-z��ʸN
���`���6j}�g�mP�,�sF�S.��C�Wr{�� ^`��Q`��*��,���S�q�|
��W�P��V
9g�T������r��	�xzC��aZ�3�����T�I�P/����s��(2�+�"9�Sa�nյ�V��j���h,v]2tK`��r��mi�͸Q��|��E?BbKH@R�.w���MHOA|�1ŉ�&�1�b�#_'�����+N�^3�y2�>!���MȺb�Y����fY��۔�f��|�l��=�QQ�so���'L>bq�&z�>�i!@,�R�x9x��%��!#��j��i<2���M��2>��QtAƘ�|Š�m�_B���fH������j]i:���\B��-�=�$	��ו@��d7�q�N���Ɲ�p ���S'���9k�1s��k�}f��Л߃ �2~�i�u��T]ofED���a�g/�`W�X��xEk�e?�i��`�i���w�\4]c�����tfO�6�
U����_-RO�dam�����F��2b'��Q�ح�5�hO��v���bMbM���%2	�?��@F8�QjUDU��D�m]Jr1��q�}�z<�y�?	��v9'�${�-���o�T�_Dt��ܺ��kA�>]rU�5��)��߇S$2�W��Cg�Ő��uu�4�:>�
���,�W۝}���pۀvI����d��8?������a�NL`0?��u����s�M���i��U�gH/;����0�u:x�g]-��QfR&Tr�J�̞�����ȯ^n���v�Y��?{
��/�������YV--�aP05�0ܝ���J���&�<�B���Q�T�rrS&���j!4�G\���@RZ�){���/�VG\�?��'�I�r�������&g�n�����2lY��\�p[ct�g�b�~���J?%> 9��E7W�+���ƍ$�(-��Q�ԏK�r3r����->Op�N���`tO�H��&n�ڽN/�k�����=��Q!�Ie}QԀ4g�|���95�
'	J_�P蹩���4>�X� �ݵm��T2WwD�C#�%�=ڼYST�C������1�^յ|T�W���������ʼ+tm�PDu�a�O�I�*�:fP6�)���E�V�F��S�Sk�1�����zm����dm:nW�&��b����Ġ�tT<�����"]&:���,��-��b�E�8w��_��")�f�d_y�j�ja�I�W���B������`�?��brI��I�Z�t����c�v��a�8РW~��j��=��1�j/d�
b��rp��Ϋի���$i���u������i|�u��d�#?��I�r��k�iL�ۄH�r���N��*s��F�����Z�J!r��1Cƣ��-�c��p���&��Th���eȥ|)Ȭҵ��O!s'�K��x���F�dᶶY+9��[>z�aDے�b���ȝ�a�bMdm�BX�c���\�"\�`U�����>�$��Gp|3A��.���3����Q;��*b���E �0��3��p������>轧 [�i����a�A�������7F5�������,1+ӟ *袳�=����~�?g��VC�"�Ȉ|_�/��mR����&g�x�p�"���ɞ��ّ�!�pL�T��a7����`8����jU�+�촙 �</D�u�;��ES=�$��z/*VL��JG�jbⴘ�C)��V�V�=��|��Ѩ�TJ"'��XF7���I��~)ҿ2���tE����������!����A&��x�"�>��h[��IV�5�� �ѻO�V�Q��6���c_+*�b�>z��7�u�P̬�\��x^8��&|�0# ����T�ʋK�E{�j~�!�X�=�^ %��! ��Bd��p}��[Hlb��@��_l\�Y�������vWO-+n�Fǂ8����E�G+V�BN��r܏�<�a�{��R�
���1,	�Ǳ�Eu2�hw�Rct1��^�};}[��?+퐤�\6Pl�Hl�����g���<CȖVI1ץB�Y$>�b�)ȇ�J,�MbZc|\,��7z\R��^����nѻ��r\ܢ��L%xW�J�Ƚ�W��2S��9��j/8���X�� ݙ�?����d� :��p�?@v���{�+�U,���q3W������B�?A`�����e�ڌV�#��
O��iU��ȳ㠴Zn�:��	��L��`}����+*`�F�Ѣs�nPng��n�zۯ�����=P)~a�s���Of��l(d���tV���1-�LԢ`�����-Qn�n�	��N��B�PW9�T�1"���p���ip�D�p��Z��]@|�+H:��;&�7Ja�8����X6��Fs�ߟ��y�E��,ĖEY���W#�5�K��o��ۤ��
���Ғ�u�R-5g��:�8�o~��L��^�yL��B���8 U62;GSy!�`�ȋ�:��$��
�ƃ�r8�p�B���󶤮<聂���a��q9q�X
�O47;��)?e��w�^�O�����ֽ �>��������I�OS<S^������1v3}I�9#ݫi�#��ȅ��4�z\���.6�8�����Qv�^M�I��8.Η6��D'�>�j����Q!4K!�8,2df���ȷ�Um]Y ��R6D�7�wqO�}t��C�(m&q�^�K^tYۙNLv=J�P� ���% ��\��� 칚"���W����d(˗�|�D˓��9a�z�Vd\���2P6���k[A�5�O��%�8/�(^�uR���;|ŷW怅.�����Rp��B��Q�JR{b���v�V"�u�/��i>�nLAص�S�s���H%\Hgo���t񜂧�91�[m�'&�E�w���T�Bp���mЀ4�w8�2��-��f�����Y.R5���]XO��+�^�`I�ese%X�^L�^� "�$e�*�sٯ�C��C� ��~%�X${�0�6�4	J���`�n�k�����t��T�Wj{a3X�+q�bhMS5�r7�J%��̇���ot��'ᚺ1�uۻׂ��+JO/�\*��)��*	t��P@���K~l�~2���2to_Z^5�z�)�{"k�����}�����:�R^�'�8)���x9��2D顷�(8�����6~���%��Ǣ r�t z�U:	���D�C@��ޖ�g���U&v�;��7f���6��H�
�F�c�y�w���K�c�����poL�h��%,B��F����q�-t�2��@~KͿ�Ok��@)�\-�%�5�e'�1�T��P�z@D�QR଎W`s��	�nXC��.R���!x��n�6ij̗�	\tx����"�<g�-�����`��5�Q��<�MgAn��˖:��T� џ�whC��Abo$�`u�bv�f�}&�{�݊��Q+�]U����Ѝ�	���j�<��g�m�c�͂�;}��i�T��:G�y�ͪ!��i�_pc�>�L��9��PB�A�J
�r���Z�Qo�!�Y��h�����Sf���a*b��	L��n��z�U|m�5/2�c1%I1]���"������1�K����l\U����X~���ݜ�fH!�Ts��K�!�*���A����l��
�V~a=�	ʝE�o��^����]r_C��
��s���7l��6��jo�E���;�Õ�����[��'ɯe���
��i���<�Nh���S��Σg!|��:�`nZ������~<�oAF���E�e��ӭwZ+�j��%J�|<V��ύ/,$	=�%��>��q)3� TX��If5�$�m^�{Z���z׻x�QrqQLM��H�o�@J�g�,�����kJh���Rr�u)�~�J�CLI�����c�� Y�3�g�������y7i��
,�L�2n�F�
p�a�y>�D��mq���@����8~�ӥRH������05��&Xzf�E���>��ݑ!���7�#�8(Z�9�M�1��@�q�[���L���]EH:$J@"�L�����LG�jt_�P	�`�}��iѐ���ܑ�u�L9÷�8JKWĺ�U����aK�?��g�@$���p�<jNW�K4Ցb�O�A���'0�6&4�WLt�P<���A�5��i����'�oS�K�|4��SrRˑ���;���8��.%��@��]u�,D�5U��:�E�sp��͒ӕ����K�V��a���v�d��"��Vp��i��r�5-<�.B��M�G�P��˖Cp�&�}<NǾ�dö���,'³86��i��o|�k�
��pâ���@~@�2���!�jL����L�d#������~�ƕ���qd��l�I���8�¥��
Cj?��d�b �V[��p(����g2f������*S�}^�ٴ�bו=��-CVwR{��wϮ"�sx�,�w���~k�d�u*�-.o�=���{>������B����4b,A��G�� O2"�|��Q�R���_�f;���ʪ9�D (H�M�>�H���`�$/)�vή�A����,$^ۓȘ�����l���
��/�#�����n��/3�ۅ ��Up�ȑ6ůzVhqd�)��~��L�^跄�,6��Ki���xK���u%O]� �j����d��j�7�Ŷ(�F/��A���klO7�����^��_s�k50/�U=���f�,=�7-�u����Q��ʹ�p�y`�,]��lQ0h�
���#y.�8��}Y�� ���<+U:��'�z���TD|G�:E�6{�C���#�u*���Ƙ��D��)믊 vܡ�MM�keW��Gq�;i�&�T-��AE����7h\��/���Fꏛ�Y&x��Є��;�~���a��e���PBE��R-��������2Zmd�r�2.n�c%��	>���pأ��"A�>��Wxal�������uwQ���&�sa��F�?�g�ar] (��1H; Ԉ���=�ܴFQ\�^ے�!/jB��@1�W��2��,VQSFw�r?��r�ɪ������뒛BWK�\'�t
�.@�&���=�!����@[�)��s������js���b�g��Sȉ"�R�ej|BX@e��)����F\F�gA���tos}w:Q2e�cT���nS۬�^~���Ӧ��6�l�]|s O�̆8�����o(��;]���%��;2��{�_~�
e��f�䡟m�v>���1/�װi�^D��#5r�`i��X�T�$���Rr�a�,F��%'���κ�jz�A4f���$����dr]eT��B�UX�p�W]c�q�ג�WX��ƪ�ϔ�:�+�3��5�vY^05Y:@���Hh�ę�� �k��.���`�
��۳�3XTG��̚*�	��}�L�|N`j�1���A}ϼQB��Ŭ�����h^�]8��4��^�5��Rb��a���7 ��]KAz=� �3�j>Vp��nU�ǽF�k�?����W����e9l��@���\�c�?��A�T8C:[M�OH�2��W��c>l��x��Hg�H2���O�C����������U��Ы�H[�#3�uK�˪�b�o�ظ��[��n�:!��E�ń)�,�@�&%=�H���l�A��Ո�n6�I�2�#�EIc[�t���THg	G\Y��ӏK{W�C9��j(� ]�3����}X}͚��MG�y|]M*y�+s�y���:���\
ͪˢUN��}��w��rc�h�FrW�����U{Ί����������0tpE��x�*ף���'cre���n��gz5�C	���8_c��_ �6f��f��L(�*^��7��k�qT���Ckw�����{;O.������1dl���ή$�.f������^��?E�s~Y��K�$�NxL?S�{<h�?t�D�x�_�`$��Aݔ�:G�cL�]��nI�F�$��M���\ӣ��	�X|���T����^__�Q]ď����w�h�jŚ�tFe�����ڞ�R��d�(!}������/,���I�Bt6L����h�^hʱ -֛�u"��/s�0W�at?��R]`�D�{��z�!�����uԱfh ��BH߿]���P�� l��]"�%�⃆%��J��	���h�8��8zl�X�5��+ǚ�2���3�X��oX��|����)NI���&�=���LВai�N#�(}�2���f��kiO�66�%Pj;��?�
L���9�q*+�tW0bn6�5��HGt�Xoeb?յ! ��!�����8�&�m�=�T�g�s0>�7=��W!%�ĄQ��	�"^!�w��[%�J��O���h�2<����K��<�g.b�=��;��7l}�V�GF�W��|~�S*��Li*���Q{}�26�DG�Ät(�on6}����K�c���ev��$��^[�'D�͗���O����Xf��5�8��^�b��`W�F�q6�^"���%�����iCq�g?��4v2O���}\����[d���R�f.g��f�o1�@�Ɛh��H��o�5awa~v������X� b�� �;��$��_�ʵd�UT�F�*ŉ"��2�^=~e��|n� ��jA_$�����	u�kV�1��[�ؗy8Um,$t@�>B<�{�kk���5)��i�G�x�\��'�� á6� �+&��=��Hkg������PkV�|�6G�ן�I�e�<�:��4�c�eY�DRFz4N��3J�G�uZ/丫4f6-���
h�����h���鉸�"OR[k�F�H�j�X�#v�Ns@lLd�Q���3p:����Dgt�}�I6�L�:p��j_� �0�Zkɠj�7a)�����`�C�U-��㜜��]��O�B�j(Y�"R\�3m>'�p"�Z�ͼ�l���=�\���s�����F��}��ף�0�~�9��EL�Q��Q�NZ��	 tF�ɩ�K9�:��J�5�bBV���]��&*��1�3jFsT
E��-�='	]cF�9�
.��t�[OY ����cc�h�8���U�0���S�Z�;N���#�xY�h���S�/]/Ũ1B��8;k�+i
�W��U���3��T d�p�
�� ��6��'9 ����]%2��K
�~�ډ;���}"��P��?�>��^M7i6�I�Dn��J6#n�����oR"	K�vN�^���vq>D���D��Ԯ����*��2��O��#/dS��x����x��<�W$	�����ƊˠQ�e����ҁ+H;̂���5{�4;�є)����t*�,Aӣ�_s�6�9~�TF{�h�u�y����k�����|�Wŕmv@^����S�f�R	��*���b+E��y���ȉ�V���Km�C}o�.Dx�eQ����|�B��z ��1J��@�
l鑵wxS����a:�XF8�nܘ7f���oXy\�l?�[��c�G����, ?��GY ?{���g�ד{+/t��gC| �S���(S�kQ�']}`�t*#&w�V��,ϑ^�V��k�L=�p��1g�J���d�Ɔ$K��\��m	��?I�W)�q��P#_�,m�i�s&�#��R������� �Ñ�J���3�uy<5)�1���y��Z��>����BT!w���0eC}M��{>w��H��E��]