��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w�6V�%{������6}n�Hn������b�w.gT��#��E��׊$.C�8�D�2V������r�,�4���� ���^^�����-��9�	1�Uw�Kǹfb��Lf�}:�"!�"�]���������(�'�ꃋ�ۙ��i���} [�gs-��{\<��ձ����,׸����H
�V�zk�=#��;=�z�-T���S^#�U�a9��Hl�hI([0&K�Ώ�,�̈w�#e#��^JS�@q./k&h5.��6O/p��=�n�-�iq	�@�G�	�U�f���b�5dc�1M�>VYj �S���J�Ҧ��}��!�
�|UT;��0�Y���i1F�2��2�[� J\E��I�r~�m��b#itJ��֑ۖP��^�C$��Ya�ץAB��<����>\\���:�0NK����.� ��#�w԰�E�-V8���[ũ���yg��#�S���\���3ЁU�itm_��ԉ����J���_�-����@h#����`Ãu#�;�Bߗ����;݋#��l�݄@3���M�ة��B�b3ɟ���-���)�T�3E�
ˎ�G�����く8��_���Ma�|�[� D�=-HÈ;���*^��,_b����U��#J��ET�xlb��S�@�ġn)4F �_��� ^Y:3�LC��|2�����+v�B��u!�\��L�B�
Q���qz8o��1pTl�_�ݠ>?��05���@�c�xL#�k���+��W�R����~��r�hH���q�|
s�Aop�炅�H����-h�K��G�1�k>@�
��,���:�".:;yY�K�T���G��N�L�G�E)1s���_�ʉ�<+��.|Q���'~�e5�̼7%�Eu�al������� �1:X�� ���K�F�٪NK�g��k,�Y7�R��$�[R�؃��t!�b�����%��.zr w�*��͖q�q�e �.A���
����+Rle���#���� �����9�?��sL�NJn)�j���e�W�s���J1I�_G�U5�w����h�-�^ �Wz�����.�VZ\� �X�&|~�ᴏ��Џ�&y�"�������s���x�����%��yB=;C���H�F�H�t]Xw�G�ߥ7�?�y�|*��bW@8s	EhK��Ƹ*��������(�Y>
�����3O{��U�WH��)S���*�8r_��F�@jV?
*�i�Fz5�����&],8�
�qp��BU�t�(�귲�x�[A�/vnJp�a,Lۢ�N����z��#���+7cj���]�X��m��m e[z�7l��<t��4��"^'o5�R�`����֯�ȁ��Lύ�-���p_a�T�E+�m5989���u6�� �|�+��嫑d���R'��;w��ˣn�T Es��Y�A	I�(������JI��/f�(�G��;�IU8 z-�-¶X#%����zй�\Uy����@F9a�q��^�R����#E���e]o.�?���<���%	�[3W<�U��Ҿ�1�}���}�*�[5(.��Yq�I��5���۷Uh ?��k�3qz�	E��w���}�¢V���E�·�s1���AE���p�Z!l_�"����l `&���}ݙ�"�=��A���K4�Wa�o��2]�%�l RƐ~�8�2��X>_�mhL�.v�(�&��ߵ]�h�޳��<�bU~a�� F�u�J���v��N\$":�����ء{��ý���N��2�0:��˷�G^�2�jz
+x/i��y��?"���9$�����3��%�ۃ?lƂ9�L���u$\W��|�wv�׈_GQ�1�̅���pf�`��u._PA�7��2��D�*����v"����)��Ty�M����Ļe9](pϊ��-�T�zU�:�����]����j����T���(t�M�l1��N��,.߲X�1j,��\Wt���B\q�Z0����m�4�?8�gf	�e4lv�K��4���_�O����Ü�~ڊEׅ�Qӝ�{�F\z#��A_o	5���f�%b���K���^��恾*��:�7�/ç�g�<� � L+�e�Gr�v9��IAf�vBI�$;�����7�'�)�1*P� ��Yf7�4���͙���E��OeA8�n\`x��;G؃���M^is���
��ͫp�/�Ua��ܗuR[*h��Ns�u
HG�[�©ώ_\�ٞq�;�˧��pN����:�g�ν�*`����v����,��EX��`�*r�������w�eL5htS��!�N�n�F�k6`��].i�XV>�=�p*_|����5 	$}~�Xv3��=v1�+�^�h�^YP��WXnϜ@��FsĦ9���Zm�&f�>Kn�z���������쀆W�UD����X�$��3�Hh�`�BV�؞����+vT6W��/�kD�&E�k�o��37��{M�K'᧞a�4�r��*K��h^�8;�z��ێ��I�ޥ���� � D=U�B�GR�r�����zf�r�J�~1�\�\�I?�Տ�k)#��]/{�R	x����J�2�V
D�!;m�0b�Z�k;$`a��APMrA>8!`�����Y�9�rଃ���&l�L@_e#��Ée7n"�j�[ ��*�-^K�SEy���x���ӡ6-�h�C9�5ػ��qkuG1��t�E��P�卪i��ȑ��{�o������maP+2�x�s���P�-&�*��h��-I�5�.b�j�t���wm�'(O/"Є�v��'�1$�_��t{f����b�Ů���DF�\y�9�U$�(��3��?>s�),Z�wJ������b�6��q;Dr(�����Ǌ�OY��X���4����W�l�ٺ�#�fi�s���k�k�<��z�!�QK�oA���'6Ѥ�Z�L�d0�`�F���t�O.�?3iH#>���,՗�1�}��9��2�	�>6����R�����5]b�EP��G�ե&BX�f{���d�������L�'>̈\��	���J�������]U�R�������|e����,��D�e�%��V;!#Δu��U�>�Du���� h�)5Ӆ�GhN��p�c�Wu1RY���p��L�Т�͞�������V<��h0I�4�\9b�X�YvL��(���Y��5�/�\m����ϡ�~���T�#����`Q��ݡ[W�(��#���)Z��x'G*v�����0V�R�l����3�y�Ƌ9Z?j��w+�9�v�'𭯊�C�꬚4�d*�Y�+������f=0���蠳&1e2٣�[��0�8��%I����^<)�-F]$�>����H�$2���!��0zYp�;�s6]�~�e�/=��4�(#L�����.|^�"����2}i@��Y��V'a7�*���|U7v�Λ��~��h�Ej����q��ż�Q&������R[�[�M�{�+��^�jށs�ƌO��is�g��1p�
���O;���3��y\l�����O�'L�����30����u��=+}�hr�ã�����Q\��б��@�,�D򠆂�9��}�{�d~NQHt8Nʶ�/u `Y -�<@�P��@T4c6e�����s��^S�P]��O�.!�2������eB���Iv�=�`C��.J�=��������wdC+��x- 0��'�wZcLP����8Ri��Zk�$�T+�p_� ,�5�G�׊-
� Dq�]�bZ������2���ձj�` ���l��N*O���ك��a��l��-䢄�mjh����<���?�˗|jo�:3f��%��n��[�M���n\Q��$���VU.��,6�n�(�U[�8>WQ��Z�GC9x;/�g�T��'�U�N�������?nwg��͈~�T9� (��9�0�.�c��.u6�uM����@��DCɌtZ�F1�Yћ/�y~�/j͡� <;g�LQ���e��������;����we4-yʹ���kX�|�ݹ-��c%��&���)>�S�� y�S#�&���Zqn���h�.�FEu[�U��	AE���Z^�Y��
��<���sE1\��jKt�tؒ�@#s^`}i\"UI`n��o��r(���:ѐ��θY:���.ϲ�P�q��X�B.. )�)�l�3}>��u�n���-yϬ��_�N+א����%v�}�Y�Ulu�;���� � ��إ�>��&��@��D��K�<-�l\8�P٫�Q��Q��~�`��]J��ݜ{�R��� ��A�M-j�u�sLoM �j	����D� �w#���y���A<�n�ŵ���=��wВ����oH��J�Y�/��%��L�����;K������#zP��^�6㳦�#���QCau4K%~1�n��Q�7} �9D
{^�+fi���%��Z��^�3n�RM!^�;���f.�j�+�k�-� ����W�<W��\z�S�@7���'�hTX%�Cg��b�Q��iM==A^���͙(Y*Ѽ-������� Q���Y	�s��L�k� X��̿�	Pt�IU&A�����L����qi��aF�܉�[=���U���ljp�͵����7O��Y�O��(��l%�+��q]�8�؞����3�r�7�[�h|�ƂD��v���Z�X;�f6�G�ҿ��4�z�e[ G�w��bv\ .HL��Sgi����,s��m����_����W���$��� �}M��T���B>����o��C�������]GsZbOU��y&��*|ث�Y�
�����y�T�G�['-��#6��/Q&�@w����_ҁ�HU�:9�Xn8I�
�Ctg��V��^k�i��8����3�ǔ������h�m�����hR&��[�$BE�jm)r�^�ۻ�9m�1Kב����~�-� $�?*�`�9o����	��ګa��c��`Ki����:nC���K<��?�5S�$��ټ�����qj�)��Er �X�?i�<S��t�D�)�&S�0�D�q�,Rc�!�mR��B�q��wx'E@�m����U��1X�{:"��}�q}��C��iᖩ������A�Zuub/��׷��tgǱ@&���� 3���}
�Z�`�P&�ѹ��nԿ��xh��v����sZ���}gM���ߙ�*E��9�'��`�cƧ֐z4��o��&o�ZZP*�Q��hV�!}�3�*�fm�M�'�m�s��Ǖo_�U��{L_X8�+<�����K󶪯�k�!�"����i�0N��1R3�e�^��Q� �@7��eڕ�izv�[�z���(��|��Z��D^�P�:ʰ�����Ч�����T3�12�8'�d�.db�ʤ�5{A����AJ�3#׿еy�J��x%�_mdY?=� ���+gw&��]Uo�_�ѣ�V�+�x����
-�X|�m�L�-��y7Pi��A7<��-I]AEǻO��=� ��ή����߉;���LBMXZ*ˣ�v�xvS���b�0M>�h�U�<6�f�:�.��'ל��kk�����g�Ց/HB���̾����0?x��(�of����W	K��ʶr��V��=�ovsK�O1�M�n`5:#͸�_i�clPѢ;r�:q�Խv���ʼ��f��j1��N�zD4�i�F�1��H+@��hM����a�1�6u)s���މ����¿�9�l��C	>�!����"ڨ�mKRVl4n�d�O㻀�ҽ�?Ļ9��ǄO����̤���K�D�����Z�A��������H9�翲k�H`涳�#�>�Me.�YSrZܰw�Nw� bB�{��� �ߓP�a�z�1i�A�A?����A"��z�:���Հ�'���0>��A�L\�ɯ+����v��E�ߍ#(yI.㧎>pL�4=>J�b������Wx�,k^��Y0��Wg�� �o9>j)/4�$�d"��-��]�H ��y�E�"s�VM/B�'+ww/�K#G��w���h��ݜ��g<C(o�XsL?��#ẃ��yWY)��G�l9\�$�O��)��k� Ȟ�;�B��
�C	�g�"�:p�D�����o��1M�A@p:q �Zȱ;���x}����6��?Z��L���C��J��#�$SP�(W���19��QX�Vs��*m�N_�}K��}�����Y��C�C��:�PoW���kZ��4`5.fel�4��/H7ꎢ��0!�9%� DpǙ�]�c.��ͺ�VĞu�k����Β"�x�g�'.�A�%օ�yösV�#����vy������oc��?$<T��V���(m�s~���f_������y�0�\_��Ie+JD�͵d�1�'(�����K���l�?=A��;�V��qy#��E���N���KA��`LJ�͵!�d�����n>�JQx�����?#�� *Ю+1YN��s@�}nd���F��hEf���*O�'�����uvbe�0T����_/SzNq>Bh���Ӓ�R����)��0^l<m�%ܺSQQoD޲cD�ɗ`�caXA
�}�����K#Vw����=a���t����x�1�hޤ�"�S�9ZF��/�z��JGh���i��l�`^s��;Q�Uݒng��J;�e�Hh:<8C*GN1�Jw"��*��-�6g�C�Wɞ�1D�����JK��{{��jC�Wi���󜓁L1"c���a�O+*���.\�Y�^�Xn���L͇�Ց��%�fA�(�=zhjW ��S���#Ē;Ρ�� ��r͙ $J�*��vh<<܌z��!���M�
���d�����5�Z5FiTp�i�9sl�l�x/�]!Њ��+�u���SHV���o��6����r/�V��ދ�<,�<�̾�/��r/������oA��G�MDgM��mA�zx��E�Y.�x��9�V�{t�<�YV�A��2��wNq�m�y���D �'(��ָvP<=���v&��`�j V��=BB,c��8�GQ�,�{�O@	�H�64��q=�q^vȁeq��G�di�K���Y)ȈLgLf{$j���_�S�f�z��=7fe�
՟��ر��t!������5�[��Dw�
P�;���Yj	HL8*j.�Q���~��Y�N;��]�	)�z�:h;���8���@�m��#a�/�]��~���@��o��ඒۮI���7��1I�AjJ�2�T�=�X�N]?@>2�M�,����Pd*��b[$�����������# j���;q��+������# ?���S6)8W<ܚ�zإ	��έHe�WKgQ6��ϰ�����f�F%[iY��H{�AW����c��JeF~���U�ޢ��7g!�m~+<7繫=�H��h
#4Vd����%��zT
Rז�,�93D5��Χ}��1Z�I�ؐ 7u���.1�*�"Y:���՞����1�.�c�h\,������q�ƸT��:��)xg���r��G'~�	�����K������)�V��/�PK>�n�^b|��F������&��q|�
��8��4�K�����q�Ẁ��F��kz}�gW	<��X�͖�SD�[b�Gw�<΄�`�8D��n��ӈ^��&h���U2�.�JK�(�?k�����rY���|���q�}ʤȃ�4���	�V�`��8>T�U���IH���L�˛m���1n��c�l��i���zK���)��\�u��1c��(�a~kq��U��+W�OM�nw��)O�Mn@[!4�O�����#p�.Y%%\�Ak�x�����'%��`���h�1�0F��u 
��kM�
������l�&%5s��E�M�-<�Ødݚ*-v'ૂ>K�{բ�bs��?��C'�y*;U�⌹� ��	U���B��	R$!�.?��*]�"�w�n�A�%�'�ܓ	ʮ6�q�D�wÞ�$�I�YJ��~�_�]������63�ӏ��S�e[���l͒���<�~�݁�3�N-�W����*��S���Epˍ�hd�Hr���?I��7����d*
lj���\�0;5�S�5�B-����y��޿H@��q�ϾOC�����OMm�W�M���6\��j��*�K�I2��IP�hzp�2�����TP�NUP�s��J"��V���\�+˥��8��uf��������o��	c�^ �XCq'zW0uB p���|2�O����A�J��"����7S=���i��E�ʚl2"�"h0%� ���A�^�� ;���6�`Os���_�
���l��r�.6�:�t��j�E������XImm�_��6U���TOgO��n~_��`su��P�rY�����
5�ETP�����4��7�r�����T�xx�&�z^�Y�ٸZŞ�R$�fW��/�K�(���k9�2J��\>�XI{w⌽m��H���ާ��a"`'��Q����έ�{����P���m.Il=w�f}��pR`�@�` �B�Ub�t�<sR7R`��>Ԑ ��*����i]��	��*<�*=�x�R@%��լ��V�9���m��x�����k�|V%"�2�Y�ng�?r�>n �<9���w[������"´̲��[&��p���%�Z���>v/c%���37Mv�._��q(� Ւ��m����޴��H"���_��&�p�@?3���2C"����ϊ)>�M�;�:(���[�d�A#��wd-���S�{v��ލ+���9rw���(ޯ.5}�����_�����xO��B�3�mh��ƣm��?�;�]�$�h{T��+�F�7��,(���ل�b���t��3�>�~6�&��9(-Fj= '��NT�4�~\r�7�h�(nya�W@4See�f�D2���V�u����	YI��@�
�������%wQS�ԺUb���~d�a������t���ѳ��NE`�V�抋O�j��ګ��}l�TG	�0Whs���
���֗BbL�Lp���{��%	��\M1��$E�#왎�o�ҩ4�ˇ��@3��)�������͐G	Lf�yVVњ5=�.@O�p�c�_��^h�j_*��j�����@8��}�vE W4�o9u��U���B�_���2��\�Dqm(7w]/�_^��j�y:A/%��~�~	>�f쥿��rв�Ec-�v�� G4���Ҁ�8{?�UjP��-�,eU�����+mQ/;�Qb����ﬀ�Mt�_��=y�c���{��v	W�+s��o�Y���ǔr�k{Ǖa�/��l��H�+8��^ef��'-�- ��ݶ����<��(Q�7Q��N��q�7u�J<0�;��2�3�eeq��b�>�����3"��H���9�>�6����_"do`*3�������ېѯD�!�[�Px��u�?���}:܍�0�eu*��R�;�
5�5��	3Z����qr��R�Z�#'](��T0a���pAVU�E����� ��e<�^"���m����句%�G��"_�_=��q;�D1�)�J� r�����ʈ)�����
=�y�p����O ����(���4�"dc���XP�8�A���h+�9�R���e�ӊ`��¡�*q���2(�G��O��89�Jټn9`�Jk;���$(hR�6��@�,��.�"V��7~�vN<[�M�h�����d�3I挃��Cz�S" ʳLK��,si�Z�0bL,F_��l�8>���Su�Y����YΏ�k��v��ԩ}��W��%��S�Ϲ�E6���<�X���G(J�^�"��3?ovm�u���+6I���j��/�o��q��ғ`���GW�m��$�%s�i���	�F����(ٞ9HKR�Z���4;�	��Xo�a�0}kqr樋�n��4/�i5mʷ��YY�v����{��@�zE�$!�]9�k]mw8�� w:W�\��0I6���pS��b�oY����!sL�ș�Nt�|�XvO�yx�gBR���Ւ���)tW-Dd�'�2B*0/q�Q QQn�A�u���g���=�~��9۴�X,��K|����@#ֽ
���_��9)۹����Dd.2o��N�9�WG^3��3���	���Lj�2V����v�M�"nt�GP��e$з��9k���� 	>����g� G	, ^?��٬����[o��8Pi&��6.^��BkR�Y�����
h��S�<h�X�	u��,p{���~��	����d�����1#4��2�|9 �Ιg�;&��/��� uW���3���ç��8�O(����T�'`ᬇ�-��~��1-^]����=�

KN[�����X�:��B�e�����j�N;�W�Vό��3�Q&���+K�㿂D�����S\�s.U��5�-�тL�1s�R�(sV�	�"�«q��R����P���y��>�8�z/t����P#�ԋ�rZ �OJ*�)�Ԟ��_�(ǵ�(Y�]����.^qQ��6 �X����$�{��ӕ�G���T�9����i@!8��"M�T�"����V�^})�xGυ���R��+q5d�m�`�PI#�я"�ٶ�[�,��GjT0��a�"Yjۯ�aư�qF{��x��+�{[�ͳ��R�$e��F�lᷓOL¸_A�v�U�>��N���ߨ�[% �eպ�;Aj'����G5őe�?L1{��@������]���C}ٖ���W67�M�5W*IG�>O�Eֆ)jS��ﭷ劼��[�������ܤIb}��
�u�|�ёE�f<�?.O�u~�3&�$ïkT<��։��؆ي�F(�_o�,r�����ѦV���@�d���Z�����e����j$�-�q>~4G�j��ͷ����}��A1�p;)8pe�	��ɜ��&aZ�����W">�o�W��J7��_< �}��Mº�If�1�%��ه�J�ʈ��.��հ/�j�������Z�;<� �J�������j�>Ngz:��(��^~��/i�2�2\Uc��J��B���onSom������4�㝟HH��E�V}ف�	_�2r{������p8V.=����d�f��ܼ)���O\2o,fѵ^�b��9�
%N�#U�a-M�ހb�z�2ԉS�����+ӠH�
i���Q����|�I���Xj�cgp�VJz'
�
gJ�l�؇�7:�L�u8��0ڌ�2�H0��G4�E.��q�B���Vŷ��d"ߚ�/����\Xx��N3���!SC�AZꎪkA�<M���`w	��f�!X$�ڄ���R�[<���5�qRl��@��ObN����J/�]�\��>��<'�p����wM��a��F�r���%�-2R�أN +��B�K˫T��O�g�U��`�6�v�VqhvU���������G���QI�$5��=O�w�5~��y:T��A�#����J-r�jL���@�2G��Z�S�Q0�]4��x#$ԌkŠj~C�Ɵt&0��O�U�}��s�)g��GJ�s�nR�P�?V��'��xH��-���`���:/��J���ҽ�@�K��,�^ ��*���I�|���0��r��8�"����s��{8��}��t#j���<��)>K���k�Lr �%j�f�A����{��"��"[��_wAt�n?�me�̼����5��c'�d����L�v�ER���U�u��Zض�K�?D�ΈK+��v�G����x8�ޜ��6�����!�^��"�����B��eY-���{�#7Ƞ�,��7�ն�'��RI��5������P��O{`/Z�7��%��
���1�����i�H ��?���&���
�Rׂ��E�>�v�r��,~���r��K�����LM� ;�H�����/��H��l%t�7ߠ�B�v0K�8��}<a]r4��_BWXB��R v��J]�Wr�r�����i���B{ƕA��>�j&d��O�7B��6�Hrf�zq������{�n�k��U�`\���cm������U����Zh9O+m/�	��h�W�X^��?��/*|gݾͶ\����	>]L���i=h�ͪ�F�zo�kD~H��9��q+�o�"M��2�i�{d2�(t�����<��C�G�?F��l��MIѭ�qMK�w� �~����l�8�}����UYx
tK�cY�!�8�u�'79�zdB�ڋ���[Bzڋ��	J,rcRћ=yQ����hW��V���KE}�o�<�S�ϖ>��C���O�R����&�M��cX)��/(;+�TB܀������,�no5vLѮ&�-��`��V�@Cb�ǀ�{�b���0w@�ۖ�VB�b�h�?�6���9� g >�]�["��;?u�C�a}�4�1)�M��ቇ�Kx����7�,���bw���Y�2�RO��Pl��`�hw��p益�����2���Ű�d��:��!�����C|wI�'�L��Z�Cd}�w9W�EG0B��a3g̥�-���:�z�C#p<	���"�Ұ�̧�l��4/ ����a��7��kEŐR���.��w*���%L�k�:����p�
j��%<�*Ձ?x���t�RM��I L�Bà�i�O�Jb
� BjQ"&���$��pJmC�η�95); L�I�IA���]̬�T��)�kI<�.�����.7�H	>����"�,��F3]��TMQԲ�5���,q%��������պk�V땴���û�<�D���d��Q���:J���=h]6t���w�T,��%>����:!�f,Ll|��dx��;�5�^�홾��n�IYWv�m�ؗ G/���Xn�:�"�PB�9,��R]r�ѥ�Xf��}9�w�cQ�,�=)a5�UڎC��W6)�D0KB�0��a<[��>�_,ƽ����=Y��C,Lؾ���$� J87��?0CG����j�J�U�kD�������	�3�?�h�[��8&�����$��;L���ʚ�a����I�+d�Υy�� ��S�i�u�TzyF�H���6��б��$�u�ݺ��Ʊ-A:��q�Ң�z�C� 囟8��Z�S�����)��*���~���\�y
����6�r�{A�g]Q�9Jx\ń��eF��	7R��s�t���DɻӪ��c�3.Į�-R-z��l�s5��G�����G�Ū��N3�Z8�N�hf>����|���V@�zm��0%���:���95��A����G.��|�z������)�C��`,����1��;#G�k��ο�b-Yl���&5]Ғf�)�a���)��!Y��:��������[=u���I~gi2�"gKc�y�V 2�侽jw��8���S՚��tw)b�`�Є������/c�u�e�C2�k,1l������Ճ�@��B�ֆ*Ȋ隤[�g�|�ɯ�-�0e�N��|��o�_����`����VSC���*�˞CQ/�&�]�ȫ��#*l�^�^�M}:�W�?�������Y6.��J�NѽjӉl؋������[Q���^���b]a<�G�#��O�ZC?1U�b��q��p\�#���|����L��>�w$�v,�?yD�+�:�HE;���m5N`��7%��%��l*��ܛ)#-�۫P ��"t���^�;)w&}F�IQ�><n9��R}���F g�,aʹ���T`J�Z����~�.ނ6�z��5��O����Q�z.擴 �ޭc�F�1�zl�p�t؋fv��~�_ϊ'�6Z�m����{djR�����\o����7����._�Yɝ�;���P�v�e=E���e�F���(���p@V;|����������P�~��Rq͙sʓ��h���Æ11Tb�p=�ptEtN�r_��=O?��}��p�W��S𺦒
�d���!��:@�Ρ�Xw�a��/������}u{hU��鋐�W�����+��clڜ������F��2��k��mXS�N�PSv�U�o_��t��*oں�9oaM6d8i�9�[��B�C�L�x���w7�� �6�b�[mi}�	�'ص�Rx�(����4�b��Ջ�����D❜���V��(�>�XdsOi�L���X�i/�G�<����{����t��y@؍i�yț��@�⏢}"�DbL&~�$�龩&�&������h���`�R!�Im�a�#� �goU(�D���d�>��"HW��X:�+Fy���g7�넎��P���9NH�|���|)y��aB�=�q$3�_�35{K��1�#�]w�Z� -kƚW�w3�u�~+�V�s���8�xڇ
��`�cOoUd=DaG��G��-	w4�/ƙ3���,ǅ���7	�c5$�k�Uv��ɏ�b�?�;��P4���FO&�mڐ�HΉ��h��9��i��) �{����� w�{
S�����7����집 ��:�т����k"ia�,����FQ�6��&��8�M��f��8�/^ya�/�5�47>Q���H��b[Ta�v���+��$�Q?��8�H4+���-7������h폁+�m�h�9�	�cWq:�^��\a�!��4/�\Vu�����	bQ6�)n�6�vP?�(�d���
�-I+3&�C�0'N�U��V�H�ŀ!<t���v��LǤ�[�n����uD�t���2��jmK=YثH��EN+�P6kie��?r��G�u�Z�	�מ���E�f�{�Z?#$���U�<5`�4�pd�鿩��c@�ߖ�jv�_�Q���q��uY=�D\���+�I~�s�Jw�;KOIhQ:Z�M�0g�y�}y����N}\f�p�?���U�r&Kݮ��U���gf����J����o%�.%Ϛ�k�܄�B�s�����S=��L���M[G�eԗ֬��0�wޯ
�Y7͚��8(O3ȄP1���5*�o�L�Ը	��=�.���) \O�"�ԴI��O���B��;7P��(F�FŻ��\���M��|�����Y���\���S��:t{�S:�.xζ,���Ѱ|v�
Z˨G���g����\�.w8V�;(e��N\!$���K���V&yq�[�t�I�����=�M*�T�`�?��|��,ڿ^����j�����u]!�)��؋��7w�"%��i�>�B��]S�&�tC?��$|2���5��B6�C���H
	��t��3�ɉ�ix��WM�M Q�LK&U�r�I�*�PA,/�3���>X>X)A �� J�?}� � �����I<�3�1��\��Q��InN� sQ%>�����M0{�Y&w��޺5�ZR���贅ʴY���7܇'�pb��a*Z���e`��f���i)a��k���7�u�MKۡ����X���I�������b�	�ͼh#�Z�ȷ�������9�1��j�T�����D�z�l���chr=��ư������t� �����|��ٝ�8t#��1��l�ߣ�>>i��^��'	��V|L���6���3y��bHhM�ů83��A�A �_�'{�vo6�X+�)3<�2��el$��j���ss�>֩}���.[�5��l/��ѹ>�ӢQo.�S�_Y"����\H2�#3�P������3���st�� ��gz��/��ҥ�.`N��-N��gk�|N��}./���9'E�J��_T�t��fPb�Z3�EB��Ғ����I�	fh��ٱh�������Y��K��=uh�^�\!J� ���BO�a���O��=�+E�]a'��h&	*L�}�R+��w�fA5H�<�Pe��f�c���w8��Fۿ���7���j.s��#����p�3�4r��0BR��7�uZU���B��va�\����ҏpCM�.R�@��&)=��ǌ�{�[J"n�j[]���G�v�v #� ��X����`���!�W�p�#" ��bo88kŗ�ڷFnr^�U���7���S��8�/[F�w�m�|z,�4AI;��#��<5�D�K�Oct+��X.Z�����C��*�x{�$���7�Z�ւ6�Gs��{l�f*������h��oUq����X=y�"{^�(��,8'�y���B���ے
HހwX��h�`'��á�O�5B�x\HnY�����H,W��f�*R�`�`���6Mܭa�.b�
�j�îe�ٌS�A���|-���+s�r�Z>@�������̜C��0Ő��.&aa�����L�ik�|B�I�XQ��J�t�Eg��4�}q+9�s�>�E��~�5.��7�*���o������0u=$b����sN�ar�r�>����P$j><����I^��δ#G!�l�8A��1x ��T��*����k� "��d��a[��4e
W�� ��׹�ɠ�7k�6_��]�[�D����x���r��)�C��&I�v�f_��C�����H��9\�ٶc5�Ii2��*�œ�1������_!.#heGZ�TNբ{&�����@��"��ˬ�2�Z��}�|��-����3���l`6��F���;�v��;��
�av��S�D���X���'�=��L����m���%���y����L��*���*ɉ���P��!�Ĥ�R�ZP/�`I�uY�a��}$�j|���-S"em�4R� �K���=DUsMW�^ċ�F=_}��H���k��� Tx�v�J�sƉ���y�zN�N��V�v�ܦ��L "M�{$��H��k[f��?nE�e*����������Z�Ştb��[��ш��� عw�@�bj�v_�9@��lƳ�v.�JG*t�I.��7�T��.1�F�mYS���`]������g&��~�|�nc�'�b Xx�"`l��"��8��z���D�ђ}��z�����"��+h�IZ��Pp���o�������W��.1v�qր���fn	*c�M���&�[uqzZ:�ANy��x�o�g��i��.�9�����q:���G���9I%�0*,i�yCGA�WGt᪠�*�.6A^6��_���Y�0#;D�&�����c���m�Ș.(��>���5b�ֽd��6��5�qF5A�(�q�s,�J5��v �Pi����uY�=$�;`:��	���c�/|�)K|�^���I��V"����d������ϣ��4�n�{/t�顰��t0BB��z�*�b[s4�v�P��j�rFxPPM�/�1��+CeA�b��R��q_�X4�-�A��7��S^/,5�j����چ�*�&*�p��-7.��W-��qO�f�JR�ŃME���N��f#���R{RJa��x�~o�5l�t��e�m�bb�@a91K��[К�-k��`��
?�o��ru_S`����1ps��6�B���x��<iNA`)L�T2�����c�E���+�
�ڧlJk��)�k���H
R[ݣ/83�����j���-��߀r����Cɡ��������W �+23��#��U2�[�~�;%�b��An���s�Ƹ+*$�ɳ�HF������"�M��=�"�f9x���QWc]�y#���	�QSj�j��L;'�U��SB��;�5���M�I��~]�T��)�٪�R�:����֘��My�z0c��
_��,< �
�D45F~*p�Mx%���~��Pzp��|�fH��������/�@�%_����[/�Dc����s���9_�(��Mذ�T+��;�#�k�b#��@�-��*�Y7�v3���,�BZw`51�'���N�]�e�E)0�j�Ve��w�+�>'+�z��2�D�=z��U�[x�G-�K[ՒfQ��?�&)$?&Dq��U7���Hj� ;�`�|A/�N^���2C�|�`�M!]��=z�<���e���Uv콂������7�C�Mz}Ur�E�E����Π���n����p�����.ٻ�d�������$UT�D��΋�V����3G?�V*��Y�����+$abn@#���k`F7~�^+�:;z���"�u6Ó�^��EOt$c~�{��Vʠ��ֆ�����IH}0%u��zf�&����Tb#
�Ĭl����K����`wH��}�a���[Z!Yv�|>8�w}��&����y.$,7�7G]B&^!]8᏷s����3�+�e|��9�Q� B�g��q�����o�MȘ5�K �g�A9����E�8��{�>p�!�x�h��ܩ���M)���lέ�y�R�=�����YO5I�w��6��������-�(�������kHuꏈ�hv**�/�;t>�=��"P��1/d�\4���E=�u�E��$-;�������z9�:�dR��%i��2���8�Ӄ&�].�ۄP�UI�n4��1�ݵcY���jPp�ۏ���Ӑ.�aH���[1�i�������7�(�I��|鋫4����TD�ۧ��A�8�Q�:�ą��M�Q�C�	Q�,@�B>�J��b�#���\��R=�3
ZDO�?��!JV����<��L_��+��@ 	����IP�����Ӻ�}>�R|bo0�Ge9̊����62ƺ�t��>�	��`u�1�rw���j��'T�C�Cf��{���Ft�o�b�A��Is���mG��U)g�����V�]�G�]:���u5����[j����)������w�����h 	�0n�A�KJ5����fݗ�B�V@��z�zj�	Cp"��yu�Ow��Uxe�����d30>��K�7���l��3W�@d�q��#�vh�]tn�%x�T{6Tyܪs��N_� d�����?�*�jh�H'[�oC��C���ǩꆀX�~�K��6�C���z�q�%��ǌs��`�Ko�0Ȑ�)
�!)���Y�r������
05���{����騫�z���iOJ��.Ȋ�D��y޶&k����s+�-9,��̅;�ë��^ft�&Nm�@U��K�Ĩ�j�Ŵ���K�@��Gk����^����^�*4��Vq8eњ�[���Ć�R[�֕�f�q]����G����6z�M��?gYrO�dQ8�"!������'��D����Hx�~b�R�Z]�3��.�7��-ƿ�lj�7��Hu��7��Ea [g<�[E�[6�v�P�.zt/�N|�8N��^.Z��.�Χ��G��gr���{��c2�h���O\�0MnE�3h���B���D�~�ؒc���}����uD��z��X�̋ĭ�g�+<{�mb��RP�q�Zّ�y'��I��Byb�3���}���^�c�^�Ǌ��E|�ݢA�4�r�	me�pOy�,�$;j>�2�c�,۴&�)7~���0�Rz�+h�Wĕ�Y'[�5,h�3�H>�x���Y�����'��^�n�,����c�6k������@��R��Bl9ԥ[\��f���bR�fe��Bڰ��.h �U;@S_��z#Q=?x]P��n��m��B�_6�Ԁ���&�>���q�>�ܸ`-Jw������z�F4�p<?�J��	�7�pJ���	~1���ʉ>�8R=	�Xc�} �*ӗxfrE�M��B�~�{Q)�; \��ڑm��7���� ��2n+֐@SĒ\4��  ��S�l�Xq7y��H�a�`���TV�n�*��@�ש_���(7�*�[�'pH�N=$J���֧����<DQ_l~�R�'5B����7´�׉E��Ε��s	��K{8��m��C���$&;ܟm��[>@�ĉX�2��&�SxG�~��{2m6��;a+���T�a�iL��%�F�0�����3fo������S���+]L�	�����gB���+�8L���f,����ϭ�?�����t�m�,��\�������}T�s����]1."	D��$8Xvc,B�:���HkW��Ala;��A:�Fu�I-�
�y�i��E͞wP��!�D}V>�}��_z�(���L�����.����EE�0�:U�ۢop���5:�x�n`[�-EG���]������~>�u�͒g�5���%��u�cD�g��㡇�^lsM����{�����n�j,�N0�S�[f��8���g�]�6m^Sm��h!`S睆����躝0��{9���b7_'����aaK���/����
��������yY[5v��D�+�sO�tV:�	�Y�>�;]�lfH�#c贠E����u.�жw��e2��@>�����t��o0��YB]~�]�#��ֈ熕�O=aEq�M��J����U�r�bA�������������[ֆ)B)w�sˋf�d"#��SxE��kC����D-!����^!+b��?h��r�7����ؖm�\L�lZ��5���3��izcԆʝr��e�=�[��������QlD�e3�j+����zi�Pİرش�<��p������f{ F�7q*m@�O�u��I��ļUO��'ՉH��\�)"ۺ�|[���9��K���O�����8.NX���SuV��$Q��26��L W�鋎����Bn*�f�(%�)��^(b�t�N 7j�>�Hc���_������!��O'���Z�qr�e�y3�`$����� �� t��~=������;ț����^��CvI��{�Vp(��W#�c��D�5�;�:�@;f�8?��Y��5��=����u�p�e+S�=\h�Nlǽ��A��)�ч)�P&m_�~��71*@sF7!��j|�o</�n�?��-@���n��4p;��A�K֚�t(�����\F�*�\�A>����w�j;Z�)���� ��JX��3K���M%�
 N�A��|���L��$W�7�֬�b�^X͆#�|n+	����� 1^q��i��m" �.llJ�:�O��
�/���
<��Jg�I?�c
8�"�1��!�`;<�zww�y�9�,��6����5M�M&p�UV���,���ij�
���{�@c9_�������%֪aB�^ykU��.D+zB��ĥ�m�Hw�V�M>;�)���5�������!��?�.'P4���OX���@XF,Ik�[��p"�ƅ�_�j��g5S,���`}N6�s]֑};a�Ʋ+I��fN�vO�2�z�%D`���3��eaH��_����	k|2�rE����@!���:y���3�������-?����ʦ��b����;����@^��7Pl�vW�{�T8������?��5�_˼+�GH�?�X�	D@k��(��'��ô
�e��S��Ɵ���a̸�����!>:j�]Y�����\���N&6\���& �Ј1H0�N�`�z~Ԭ������� �{8;��X�hRL ��$i���8���*tX�v��b����k�r�<�楫���4W���U�	~��>Q>��ݦg�;�'�dއ]������^s��qBqi#Y��H��Yt�iAHĘ@;6�-��Pe �#�x��O̵�>J���fkwx���J����O�bq.����a���������G:{N	7�Y��D6=��(��y��;|,Q���/5��ȷу���B"퓏�g�-���CS/	u�����8>2XČOeU�}�z���>�������?�ۘ%��������c~|^0�/��+|�ɗgl@�N5��6�bx��Rgl�+6W�'v\@ܡ���	<�D�x����)�ݶ3��=�o9�����Xxޚ��!T��=(�ܲ�~H�	��MeSOq�$܂ӳ���2���'f�}Qj�-�ɕ�kJ�����c��=�_>���@꺑w�?!|�h�X*�^R����u_D�cJ����>�Y��Gܲ�r�Fũ2��`�"����t�#˖v�򑴺��Bmk0�/��s9r��*G���t��,@MnQ�G,�C�E������%61$/�0 Ď̓��{�I��p�G�T����P��ØvL��I2:� s�f�v3���Y�����5�J$��a�2�ˁۯ8����5�z`(*~���[�}OD�.{��6���T���(U�h�H�����\?K���~Z���X��g�i�[&�
u̾��@4?��م��FY8|�S��/9��#�ؗ`�3�)a��}=6$y� �$'��#��'p�i9�։�+�<��@3 {yCQ����Xe���є��ֆ ��o.U�*�.�>��� �)�=d�^Eݫ��?��#��7ut�@�{�3\bM�q�|�����Z*��%���pϥ�n(������k~uƊ������F�'e��TP�K��#C��M4�TI8v�|m|���V��2P�Z4�sɷx����*�ꮉ"w����%{N��SK";Hc� 0�����S��K���c�ܣّ��K,k����s�����f�� �-�yS~�A���N�LO\'!��E�"�&Vͤ�d�����s-���tn�T0K��L�NJ� ��Q�w��.$y�Ⱥ4�����hl�͙�:��A���.�Jpu��G�����@Vq$zӑ��I�}5��4�o%\��W�eH�f��OX�*�zzl�
����.�6o��������JYBd1v_�s���T��
J��W<�CЏ}�8�Ύ�e ��z�X髏s"U���w(���&�T��VC�}NfI�,P�) ���[C/��nH�7x+ܮ�Ŝ; �G�7�Gk�7 ��U(X�Bh���'A��7��
�;
XV7�^�M*�&5�B�\����!ȇ)m�)�s��8���Q櫓+>���K�(�+�/�M�X�㩳+��D¤̰rh�[k޹N�GM��,_-�o�]������cMn��?;��|�6ɺ���
d�7)��}V��W\�.-+S�!�|���v𳔨� |M�/4N)�47V���r�\��"@�w���tT��W��̅�`���Ti'U~_��S�r*4�X|�h�M�]���8�k��X~��q�W��KD��*W/o=.�>������z$����I�:w��<�D��u'av孒g	�Nbrº �ڢ%3�<����a�s_&�{�߆:�o��M��]���~H���-<��ST�+��|��Z�k��<m�*���{��&hQ��ɔ�FH)����U_[.k{��áh^o�ia�m��SJ�%�~Ǟ���ݡ�g��D���[o)���5�G�7*��D��B���m ���H�p9I��9Nm]�v�P�Qk�#��u�6���ͬ��2�-G[����2X.��t�YL�t�፪�J