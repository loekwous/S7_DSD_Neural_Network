��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n��WȥrP�����S�Ք: *��rc���o���YLc�YC�O��p�@[䒑���G?�s@Ge��T�oz�r9�'���y&N�`[�;�` Ն<����t�.�Fi���D�Qû����!�}i��c��]�}��+xxցt�'ng���c��;��6g���Y*��ı���"(�t8���)�$D˹���m.���~�����;<YB��5�%�ba���P����g�D羵�d���o8���a�� ��Bo�6��~�+����4g�AHu	\Lw��1 ���_��CS�eI7L�|�F<���n�xs(y��"�G��
��_�\^	n��.&[Y�2M}u�͐�Z����f��9W&�iq�����g��掖�CFOܭ}���/����\� �g��,z@%2P�b)_���L��H���SPd�=����6Yo��W�ٺ���7�8���?�O��a4.d�+J�^r)[�.���GY���0d/[���[(z#䢣���L:&���ƿNg�g1Φ�L�
��f�ݑ��5���|U=O����L��TA�	��5� aN��d��6+*>?�,�R��%���q�)
��I��p�G-C��ӊa����ʵ����Λ`���]���w~hjS�
�N�<�9M��U�,ѧ7k���j�ֶ�m��փ<�b����ˣ��]8�\7r=|.�1N�*cj�;��1]H���}�/XP�(h���&Q(����N���BeUO�JIW�Ђ_ Ÿ��L=:���5�v�]�S���7�Ƴ��#Ю��ܭa?I��I�!dK`U��t��.~�M)Fɕ�)i�jGƭ��.���X�C��!��#Jj�/�}g�PsYbq}��Ɉ}�����-y���\���T�;�=y3�9iC0u�3D6��t�W���hF]��<�(}�ȸ{�!ZA��3*\�C;n��M�S0$��7�V�8�V�-!��N�Kj�����K���L3�����u�ȴ4J��m��?��dM�MWǦڒ���>Sg��PІh�������.E��yt?�W9�$`4m�C��hL	aDk���_RRH*�ྜ
,	�<�Ew�[��&N�P�B��e��+����U��]>��&�~8t<�r`���S�8��PE����?�s:A�-� \�b4W�+a&R�#_Q_�	�5���{v���mq���*�>������(�C�I.�=�-��Ed�~��3���t�I��໓pt�����Q����_��r����P�?�!���������kp��e�(�y��|1��[�C#tG�شR�1��l���zs>f�����|Y�&c]��F~�x|�.�8��ﰗ;��&��	
����/�G�0��0��l���Z�Y;�b[�۩��Đ��)6��ga��(�g؆���΁z�}��*;�H��*Ԓ���@t�%GBJ�G���~��U��g�v��`s�mʸ�0P�O�-@�T�mn6|ҟ^��*.����T*oT�*8�)gB�k#���-�~�r�~�tG�O+���+XwT[r�
��x`~�N6
0{�8�dz�9�����H�P���F�S���ק�vw�ң��������/���`���<�ֽ�+Z��Ī�-s�w`6b_��ߜ��2�ܗH~(�sH�6�N��c��(^3x಑�ˇ�1[�� �a�,�9�%MÊ��4�u��j�+�!g���L(?��@�(�8�[����]�5݄������F�3�|�*����ՍV�%�bC>+7��)I�$tޮ\���}��A����jT-	'rT�.��2Wv���j�V��~����	�	�&���$1�{,�2�A��ʴt�Q�6�x�P�E���g��=$��P�1�xÎR�YY�,�fz"����C�3���*�� �]��G1�(�e�E�M�ɉ��q1�b��{*j��p���<׈$ٌpN��+��'�����p���X�R �0E8(2���-�&��K�N�/E�4̖[b��#�em�=�)��j��*�(�)^NN�I�4 uF��h��Gőp�Wp��1RȂo� �3P���g�Rc���2ܒ�w��|hձU���*&Rٗ"P(C�����m�چ�X�KB��et�Y'�v{�
��nuDЏ�H�oO'�e��-�������U����t�j(E��)v~�Mv�
e$l�Igl��c�3=�x�]Y�]� ����4�W�]�[-=��0�{{N��4xd6�է�)�5�i��:!u���ˣd�,[w+�0��_ ��957�bLgk��������2LwfW{X���]��3��LT<��i�#��w3�#�u3��O��c�$�et?ǷƣL^�̦�B��0:�1O7o��G�h�0b2��(:yt9��:��a�7\P���BE��&�k���'fT��.���:i��A1�b�Մ-Ѯ�	�:��2y�˷�,�5cA���eܧ|I<&L%t���	c$r0 Ҳ4��Axm(�k@~i��������;������=��6� �U�X!��x�y�~Y��IicB7PK���i��L!���ƙk ~�Z�kj���LQ H��0y:-�:�z�$����`Da}�u������2zM�
(}b���\��K�(fO�V_
�[H��*_�����W��-fm(9��Z^�V�N�.� ��������yZ��b�����:`<���?(}��zDH0S_��ڍ��f��d�'�vxp����3��W��XgM�������)M����L�f�^
�TN���3�0s�� �!�QD?u�͚2��#ι9�b}_q �L�ģ\H*��M'y�׻E�6�K�֑�\쾷%�t�tM���x�ق�*u������>���Z1�	� ���Y`�NTz.?ǆ|�!�e�c�S]8�j��Y��|�����.kRn��1̀��m�._J�ڦE�z�Ո̞�`G�W�--E,Ǿ{��������6/��UB4L�nvX�m&{i$*��mA;��rj�ѼC�D������k��_�l��<�cG嶖O��$�^/�P����jИa�D߸���q� �S�2������=K)��y�� ��?�鈴�l������V�)��^��P�S|qӤ�F&�< �=,�	#��Y-�ZV����(E�By�/
��T���5�0!�ɨvj���e�_/OI�{4��B�P��!��s�A	�b�C�t��	�u9t�ݍvJ�T��,�;�[C��ي�X���]���9���}��ߚ�W���8f��T�c��[P ?�`m�(��%�#N�j�a���
3��t��%�ǐ�ѯ����'�&�Au��d�-@^��E�7184����!�d���#tm���o�4�O��a��hO���>��].�&�b��\N?D;S�=�H1�&��Ρ�('���r��!3�2� ��Nv�����vt���
;-�E�/�c�M����'NS�*���Iz�CDsCi���KX0�FM�^�G@>��z�@3.�9�a�ߔN� F[��g�o ��m t�Q03l�2��Xd���mS��`+�խ��&LUQ�{�#����v�%r�x�x���h�٪�_y�����e�w�8��m�P����֬QS�=��6!���5��wi�5�JU�;]5��@o�b���S�OZ�e�Y�	S#���!�-s����o����VR�-p�G��z]S�:��7/,�<^�Z�֣:c���[
�L6-�mƷTOfeF��1���>~���|���z���V��v�!�U����E\_���0�8q!��\^T��ӯ%�[R��˲<��U�2��Aډ3�}���t�:k�N�͊��R����ݾS�[����3Gc�K����=J�dP��m4�Y)�i`#�l��3,f���K�O�}h��m��o�6={N�x�����*��CP�o���bbg�e�~i`/,�s;͊��&{�O����'���8c�G%��ç�h{|�8�O�W��2��Ē��Ӯ]���	y�'���`��� ��!���#J��l+ٰ��xl@��t�D�D���A7���&��o����m�|�0�kr��Y���/G���+�]e���&f����pk18��-�xZ�!Ku������.��dw��ݤ��)�ubmrm��oq�j���,ڭ\Hno�6c�t�O	�=t�:j3Ւ��S9���K��OVU���)Ʒ��R&��]��g۶�4�5�����ƾ�M���e�3�ϲ�|�|�jF��sE��D8����B�n�bx������ʚ�e}k-ϱp�0sm~���-���'�r�`�������A!�#|�"�^9��<鼟�;�n�������X�����H�$1�{]1ٹ�m�0�'8h��1�*���g�� Y<z5���+��Q|1��!�R��9��!sy� �t	u'�צ�=[��^`:�ڤ��vԪ�G��LõG��=v�������q_����̕�#�<��� ɯ�B��}�x+�d�y��b.�m#-���(��ܽ> �^���c�q���<��_.�׮����+�l<㛾�j~I�R��/����;�IE��L쨏��g�hݾ���� ;Q��K�/���6�@uv���Z��e#ؚ�1��NUR���>�Ѳ�x
R[+X#cYz��i���z�a�����`���覿��4)��2u4��.�����tds�T'�4zH-%����Z��z���>����ru�}Sjb��Q�Z��#��֓���%xO���OO_�Q��A�Z�1�c@IM �Y���N��q>|�����Uf5��Lӝ:s���=�X\�L65����	u��f�x⏣��/��N���p�鯱��K��ZO�QO��� ޤ�!E1��</�a0"�����鲕&�X�ly�$L5�\������V���o| ��s�6��a�O�]U�c:��x�}�G�~3I��u�H�����˝��wЙ�:xI3f�-K�����d�0���f��lg���9���d���8`e�j}��`Y���v�$�l�pT��s1��S8 ����yIa9����)ZJ�����޲�^��ZzVrm�{�D��b��k7�>���f��*S������i��SM,Mˀ'em�XD�X�7�4���p�Ƚz�ҖӾ���{����f��DV��l]v�*ųq\_�WU|Z����8�\�"Z�0c�Ib��3���i��y"x�G��d�ؾZ�@�x%�c#�?�Lt�t4,W�V�ɫ)p�5���O����ح��뭍|6{���U~�N!�bI��QF�\��)F��o>�,`��"aF-J�iA �Xk���1���-�np��>��
3�n.�#'���.z;+���
v��E�`�.f4�b��>1r����M´���)PY>�oj�4��C�V1��ƛ�\+�ˎ����4'�3�x�쪒�|[O�>�-%��S��[D�r��.�YbZ�J-�	``�lb�S�L��$�D��b�d�����F�[�0��<VP`S�W]�_]|��mJhGg瓅����Mp�Ō;�n�����{��I���Zr�b>��]�3p����n���K雭�%�a�e�+mk�ʁ�%f��GI���Dfo�d���o�9���|B��s��w?�+�T��)M�8����C��T�FPv�)܎#�h��-�	z{'$C�s�Kw�I� ~^e�L#S�&�f쉌r�Y^�eky�W�P e�UB��w���<ѱ��@Ј�����%�G��V �wk>}��s�,{6���H�����1~ �vGE
""8D

�� ��+Bil;��V��|�T��RS&��/R����溘F���1����ת���#�p��p�>�
r>/�7g����0�F��g��.�1� ۨ�:�v�i
	*D����L-?J�݋�j9�06�β~���T%��e�;�����w�{�s��'�m��/�T��Q+��򪣗�e��#�}A��1|�v���`~}~͹K���G�/z[�� kF�?]����-�y�����q�+�.��UVq�ƫ�����!y$����r�LM^��bX;��(j2�&�m�RN��3�j�5��4d�Xb0����& �yn5����WM6�8�\�(���/0g��Ąw��N��6�1��uM�KSt��D4G�t��}�up+F>/�w��������B�=�H�l�N$�1L�K��`�w�{�FNI��j-�|Jv>�o��J��Ķ�Ϲ������'0�7�$�L��S1��Vac	��m�:���ZO��E�X�0sg��.�xڕ�KM6qh@�Q�
9��ū
;����C5����]C��m/����վz��S�����
�uy�!���5�T�
�L��e l(@aҥ�̺!($��c˿n<98�@$i�v��șj+�0�j�[��i�&��ʦ!B�([��N�
qC����f̠��3V2Ը��)|���aԩ���֫�.F�H=�`(7eM#	�����*#+�����P���^@Q��h��>l�������b�U�|'φD����m͙�ϒ�������K\˪�v�CE9�	�.�H�d��И]�L>3]В*1�v�J Jg�q3+�,��Ǚ������]elp�4&����]�+|B���F�%[M�# \*U�����.m.aV&?"wM���l!�J�E�	|s
��Wz��5#adO�J��0�	8K ܑDZ�ڠ��B��/��۬���P��it��ȭL���@����B圞�����Bx���i�2�aW���� y�����3^ Pl�ܐ�ʮw�}�1}���6���5"�.$���{�^�;@��Wi,�߿JTB��3z�{+j���lʏ��vÐS�@J@������>ƞ��+$l�z)w\y�bmFx��T���Hܾu,��W����Ep@��7��);�og#Q�ۥ��z8�Z���Ki�>`���q"+`��'���y����3X�������T���<�aT|w���<�r+W�)ȁb�w_P��D��k�.&����z�o9�W��h�Dq��C�baH���0���~!��tvVNS�+q+vy��`k��GM�J`��:�w��\�_�_�]Ѝr��~�Խ���Tɋ��S���5c��$d��q.YbVX��ޜVlL�Hd�7�1G�eo�tx*Gʛ�q�U�~���w��9h���4	<��5���O�!3�?�4<�=CɅ�ۿ����.��ʉ����x�|��d�_����d׌�9��(��ݘ�,�UyTy����Ϡ�zu@��z��|�>D��(�� �%�~\�9��ڜy$:���/?8����I2��Mг�Wv]�+����%*�>�������Lh�J�����d���b!i�d]�w�0�C��7�&�NO��B��df������ڥb��
˖��js�����D|����sBZ%��9��Kѭ�@��G{�S�2�ˍ�a�Mk+�I~���
�6��>T�2��86��M�?Ø��L:\�&�����mW�� �-���iS����_(�.�n�a���̤�}\Z 	�dkP[�{8h��q+��H@�x����ʹ��̫�J8A��Gꋣ��
Jq���q+���G�T��:����Vx�?0��K5��R%�C�{ܧ�V�i��sJm%b|tR���#�ghctO\�R��2�wE��}ud�l��)'��1u��м�����BLOC�����L.�а��7H9M���\�Â`)��� ��۞%9M������t0�dI:� �0�2w�*�ʺ��{���6�X�01G��@3��P��1k���r��9Vr�TR��j�?Kq�)�y�O���6��?tU�5{���J��������Ǎ�Z*�4u�$Y&���B�8�����H]1B>M#���e&`Χ_xX�)QW>�蜨(����=�=��x_��Ӝ(��a҄�/5�G��~��m)7G�oOc.A���Z�����F�ft�G~=�(i�~sb6il����]kq {�eJi�kI]����� =���j����5ށ������W��O�j�^�P�63��y4�Ԛu�|�,ͫ;�]&�*Dp�(e�kТ_�a��"�����S�;��C��z�m�����@�Xlu��������f��U*�����Ƃ�Ѥi>~��X(�y`j�~����(/���mA&���Qyꖘ@Q��~�8�ב��!آ_�uE�%z�k�[{������F)��C&����x����{�@B*��<����sMA&�fR�Y/�鮟|�5QR�?r
9 U+#"�ap.��m9C	��)U�c��VΓ2�Vw���H����� ���UWN��'�L�s�G˖ep����о�%N�a��Z�Q����Jf+F��yA"]��w��yz���UJ���\�-��<��KWHO�V�2Ql���k<��_�@��!Z�2đ��W�)߹W��U
�j�	�F�Ұ���;��F���Ods[�Kh0ϡ��B٬�����~�>�i!E:��+ބ���8�g�E��z�E�2D����Q&�<�2�|���}�j��J���0;���'1vDL�E��3' �@��?�x��7@�AՔ�_e�w9��u|N=r
�\͆,6�ς,b�'��h��|�L�;($e���S-�V�I���A���΂��͠�ʘ�b/e\��U��$w��٦��TM�+��|�1��z��Z[C� +����E瓧�4�B��7���:���-��=��@�y�w��ZT"O=D�9�d���8G��,w��S@�r�c|�$�]p]�	���)t�Y���*M3�`���~�[���GÒ{&i�V�a�/>�3%�ф� �G�~����i����:!���<�Z; �����#��@�>�<��A�x6��W�s�;����5��zOO_���;�9\� ���>9R�?ˇc��w�_��?�	WR���і��� d"��ȗ��yp�,��z1��s�
�2����2j��N/:.W�ը�k�R\�&=X�,��Ű��]�E.��ڧ{�/GȢn��~��i���������m�n� ���8���vv��9]�a�64����?�K?�����	R��Ɓ:ߩ�4�P	S�L�l ���hn��E��h�.��=?�V����ρph�w.����sU���\�M}D�F���h	��X����[�^7)���Я��������o��46�l�g��|���p�Bw$��T@M�>���t�'Uo�eRx�H'�G��^�e�C���Va�eh|?i��h��±^����J�c�>�����tp�T��������o�~fd) ��Q�qQ�=0�p����D���gȨ��F���*�YЭ�z���a�[�C����08�w�B�p��������\&�
��sj�Q��Q���AMk�D>O��B�Ee���'Aց2���+�`nf���dEV�R�3����^ڙ���Gx=)��"sq��-Yu@n��.�k;hJ���K��7��l�]�8���>l��s��#I%�� �(n>��7�
�K@��h�&]i�@DrDI �&X�6c�(���l��s78_�X<����Y�V�W�˖�+9���Qnq�>�[!�C���t�J-�Bԩ#��oC��WCؿ��Xg����PTE����T��p'�H���-F2s�[��X1G�|��93X�<t�e����Kw����@��J����݉�vD��&+�����^H�Q��������?�2�O
Շ�������tǦ/�����&�,���~�}5küGkO��Ss_�-�E�N��ut�K#�n�8it-Yһ2M]=i)f��>���]0��_V���_�lf� �t��g:ɦ����3��;2�	��.O5�;�i��̪D�+�eQ���=���-�k��w��	0��B*iC+W��vI�ǀ���~��w /��V3@�J����ϝ�
â�:2�p��i���C�v���J�d?hA�]c��0`tG�[��!�|:^}��Xk�4��TB�a/�i�*X�OIK<���~P5�K���F!�ve��.�Y�UF��q�!����cCq�_�d�$Ϟ�$���}N�zM=mE(Db��k�����J��qM����a�2\QCG[�j��(�/	���O�t�Ύ�3;*��b���SGuΑ�,�y-�����&��@~4,�i�?�D��XYxk+D��@.����$�:2�\ԩ���e�zHM��!��y� $$j��+��I�Ka�����R��1u��������� �X��?��p�D|��n�-l�x���A��.N�^�4uQ�>�2ǘ�b���l�� �3Ff���4q�sj�V =4O��S�����㞰�t�� ���{f]�S���r�.UL�x����'
���g"{풇��B-6��ߧa@��&�c,�ƞr۫&��NRnDĝrt�̋rH�Ɏ�z�7�/�ېW%.�BI
*����=y�Pޛ���V~��T�]��{$Yډ���^@�C����Zĝ�p�+�m�a>xP��v��<��UԱO�/�LZ��&��L!<EF�+�/�KCpa0�q�͖�.�خE��=��]�(P���}���c��Aj�W��pԇ�ІCǂEI�]f���j�����*FgP_�SC�b�aǼ��kp|M�b���nmkW������1��t����C�7�K���c���%J��tz8̳�Ė��ˊ�ߠ�La�`��������M��T�J�B���ԋ��nҳ��E�����������*�	����Ä�m���J��0�aB,�Q�}�6���)��?�yLWO�|�Q�p�d4�²U�= Q3`�'��tN����]���8�WL~F�Ք��*^<XMy�)+�=�&V��<��QӤ���߽Qd�e�q;��\���%�Y K�ϋ�b��	��sԳ�Rh4����	d�5�S�V��N�Oě�v���f�|�]��Z|�lX�NΣ����4ҕ����KX2�Ju���𗽁�kȧ�^�f��ߩG������d�y�J]��*	5���e ����4�)�!0<�����'�ؓd���L$�t�(I<���HiC��^�WK_Y�_S\ڥ�b�]��.��\���{*�5[�ip-�
6c��:��NW�� �lu՟hQ�f����#��s��X�Ď<7�91-����:��t�0siR�|�?�Q�q6�<����&���<�?p�@P��!�k�Sëpϩ��*������yP��l��%�3��1�!X^�+���"I�,VEz���.�1���C����7��c���|\JMy�@�����U��#O��6.�8^F�  W��������,�_XMS�?��>��>J��r�Z�I�1�:��#(ܰ�`	�?d���q��
Ĳf����	z�	�"��@M%���&]�@�f[����Sꊨӣ�}P;��ݬ�r�W�ܷ�����'̸5b��-�5���U�l�ב1,�\KX��3C� /���U����^�������-I��̩g��lT-*�� P�T�Ю�!�wu����N��&;�8<�%ш���ۍ�D��W��꽽+H"Y�ed��p��)�zf5��#������O�C���NDS�i��P��G��lAK�}oc�˽iX�n]п5�PČ�k��Nt �,h)r!-l�K.Z�OG�4Lƶ�ϛ]���u�S�'Z��i'*�.:WY��.�4Ա���T!\gqn$�#@�N~�����<$�Bڠ�w|1dj�Rt�}��z^bWW�s���.ΠIYZ[�&��Y��97CV�de��I���}tɆeX��4`]h
��5�w�<JP�D<�ɉK<������)�R$8��X99˿�-k��j�]~���.u��U�y~����P����!���ƤlZ=YE�	��=�x@�{I1B$�U7�u�:�7�e9�'��m�����&�t'���,+�Qy���AZk�e�ϫ�l�AO�ѱ&�SK��,��<Lf�T���띂n����|��Ш��a�bؖ��V�/�P��ʽ��t�����W�׺/uB/#�$.�*���7��^���[>���p	"�*�(?�l	���� [��L_���V��b���4F�5�x�.h#=4�%}�^3��B���XS���J���V�Y��3�o����9�Rz����%;f���A�D^G�M'�^���qr� ����MH���wy�o�lk�~*D�Kr���|���\�Dp/Q��J�+�PwH�ϖ���� ��ә�v���dki~�7v�En��t��tN����Y<&�Ҕ�,m3boF�����f+
�����_8:�I��A�S��S�z!�JB�:���G _*b(_�Q�L�<&�o�l���k:�!�@6�Nʧ�(!�L>�X����a@Cn%EzCrE��	�[02�WƗp1H��h��).Z\G��ݐ�ý����s0s��TncS'�R�z����FR��r�ߞg�zᱣA�}�����j�s,Z�?K/G�o
��/My�v����N���l�G�����~�-���x�f�� �'��/=:�C|L*	{��Č���h���Z�P�N����D�9I�ut���l��O:T�&�WZ����(�,�q`G���c����g���qz��j3��y~uV��އQ@��$��ǯ֐�pIR�U��VE�-h��0�+�V�{�-�}K4�e����I+���G�M�O��#_�қ�A6B�2�|Q�s��&�tт�݆a��x�N�xs �=}W��H��v���H]\d"�B�F]�t�a1�]��P2��a�:�p2w�v	�Z�5�����>���QA���Q{p'�}ψ"���1Z��6]'����6j����=�@o��)&@�DΒ���e{$D���d��F9������oҋh���E��r��������6��'�Q��dn� �(l�ǈꚼd��O�x>8�}6�z�P���k)�gn&�B�=�M�L�f��n��'0�z��?қ������vk���=UЈ6���{�o5��9C1`VA�����.��WZ�8�|����i��H��z��?�M B�324
-܀��3�І���l���� C\��;	�lA��A��3�6b(�����~�)�ת�]ղ�R�1�1�W��~�f`W80��0�;��#F��e�4G)\y�*ч=�N>�J��4�Rp�����.
w� �DE-<gML���Ue���+��N9"��m���e��N�8E�!��F�U��ؖ7lZKr�I���&�BA|T�4����CT�tJ��>�i]R�ח���%��4�����˯y+�ǘ���r�O6���<?�I�X*�5�/��N7Ot�>�m3�PK�_c��3����)���S�7:�o�N���_l�R�O��F�$l3�~���i�l�k��������i��,(�"ʇ��s@-��}m8:T;(�)y���F�r��{��lp�ư�V�ر�OK�7��v�_ >�\+S��r����\��&6č3�߇��.�(e̶ۥ�x�R���M�G��Z�0�5�	�D&��x��֦z��'6gl��rp����q��EdH�׋Y'�j���'5��9^S�W�1뛿j����C�P��}wk/N�p!4'�n�wx~!�L4=�JA�8-�����\z"k0��M�H���.ڔȩ�mZ_T2�)�)�N��R<<n�`^�AUcK�	��;�C9�|��=���wc�H����X^�K����:5Ba���}�{����6:-E�u���PM���8rN��.G7�jEȃ�>����e(VE�\���g�;����s}K�o�"�����ŷҗ��I�;�];����d%ݶJl���������9��*#4��XQ� >>�p�,�V}ފ�UJZ=���I�AяȪ�k�z2�קq<�<�"��M���)���h���-�q����YG\�B��p����9q����"Rm��%XD.�!��}�iaz�����֕���q4p���C������UwBN��e'�e�<=����Q��kG�~��<�c��nW��{IeӒ]i�]��P1a����ͨ+Up�V�q�4�"J���L��k����q�w7Yqʚ�sDmlw�1���(�������;��]��������ꎄ ]9w��ސ�S�q\[�v�֖㼷+X�A�'j�u�'���%�����hzi>�%�0���@��Gj�
TV�w���7�|��[��@��+c�zP!!7��#�V3�ʜ'v�@�</����R/��� �8�AT��a����G�R�Mkr�d9�\�%\��I�|g:���82�� ���y0eV��?����	hm���A���T��$Z����D(�:$&p�ڱd��#P�7��*���|�W�jZ~rЅ�dS����4B1t�����x񂭾]�7W.�
��&��"^j�b'���C��Y���X�i�cD�ww���6����ʬ;�{7'��߆�<�^����xb���C?�,eF+H��*h��ñ1T��ȷ��=2�@�ܳ�g��.�r�&��k��6jyv��7֜����XbM��j�Xo}�J0�75N|��:��FV��u�����OvK��Di�D4�!�+*b�JR9.��t��$n\Q�I�B��l�v&V�������͔��B��dU[�|�B>.��8����*����vx�;P�W!Q�M��}90��}GJ�����<��>5�n���7�7�"�m| �>r1�)L'����zt;o���$	��7��y��<��]A��Y�a{Q=Jg��m+c�5׳a�볆��X�� �Nh���ʲ>v)E$�M"��F�''���li4`m��Ӓ�<�q?��h8.�}B�-Q�Xw����N�����:Z"7� ��D�b�"�[i ��*�R�'�"�R)s��+QE��N�υa��կ�������o������>� s��i _�9W���)3g<�ol��C
�2��I�ۥ��Zmc1'!�;�J��/3B7��M��4WlX���x.`��nP�:���q�1��Er�_p�u
�2"�]�����B�2V&�	:o�/��%e=	_X����ڄƈ�?���5�ޗ̀)�>b_�I���+��O�w4L�n�:���߈���/�:*����I��L�%)|�~�NȔ;]�Q�����C�����ˠܠ"��`��5l�m�GR�+$e��2h~pz�����A'��
H#W����=%��g�H���#����X��v��N���4X_��c��r	�����,v��m���qf�_�s5��ݯ�2;jnP{��$���(Ӌ\�ei���q�'�˂�_M��U}{#��2��0� p��Cϑ�����Kks�#�q�KG��t��E�u�)�&��sA��c��G��vか�N�Z���j8�6�~nf�A�����o��n�͌1FE�F��J�ʤ��)��s9�?ʠ����Q�q �(½����vs�d�̥�s[ ��J�^'����I��cAbr8/,����_b��u(4�i�����Q/�@qz�BW�ӣ-�6^���(�7��l(x-����u�� $�����tNSI/-�>a_H������Z��}��Ϡ�;�!����b��h.���QW��Jg�݄T����ta����q"a�B������_���#"x|���;*����~͟����%we7pn~�vB�ᦫ��^[�E�}���
_~�)k�{ cE�Y:�D���zR�-<��8E�r���B�!��s�����$D�,x/@�w=q�U}�[%���5����<t�3O�d��$�a��?���o���T��cu�Xc�J��Wm�FTtѭ����9�Z}�}��r	luo�px\�� �G�m��s!z�����@MA��'������$����Z�y���������ͯ-ĳ�g�̴�?!�嬌�q�s����i�/`H� i���~5L��A����]�[a��bcOqM���O��q[�3l�C9m�-4���� =l.�)^3P��Ŋ����с;"�-D�y���z#)�6f��l�������g	��Jg�qp��e�S��]Sg�Ye��!�DO�s�ߐU��mm7_���E҅~m�����7�Q�ۜ���9{�r��m�:J�I��S����$��}^��r޺�5�!����8��Xy�2�JH*)Ϭ��ůS=_��f����-$YS�PZ,ܮt��$�+���3��c�\�!�m׫}�]�:������\1�G-��-���?��X��j�щcl-�'-��Q$EB>lR��K���D���s�ȡ��nE0^�u]�g��|�N�+D�֪CX�}���0Ⴧ�d�FآP���J�>G�w0��u.w[�#B�R�r��Q7����hd2'{<�RO+NR-��p�ع"���E���4X5!Uft��%PO2.���^����m�O�,�OJ1��������)ʵ�]�:X]������aM���k!G�J�
Y|g,���CPz�*� 7ܛ麉��f�0眴�7��x�P�q<	_E����e^'�T���6e<s�����&��"�r��ig�%n50?޵�a��kޠ��mt5����}3R���{sZٛJkA���Sz��`<�Z��X���6�F"j���[�:���!�u�JZY�j��i�9+� �^��`�ڋp�UA�WuE�r˜+R;�Ζ,�j��+������y $�KT>c��E�O���w:{d,ܜ"��z�Kޱ`4o1y}+{��Il���|OG��R�������_��̍e�	�2� ��v�XeM$�\�P��*->y܄2zR�
��O�7�B���rwg���
�2��>�簯�
�;�hK"�N@=�p枷"Kط\s�N|&�����%>֧��D*�K�|���J"�� ̍u+ڣ�~���P��A,�4��D��O��h;dß����m+e�ؚ�����+�L��%���ۼ�B7�SmJ��׈(��'i��M��FA8��Y���I��{��×�'��ڇ��FX��a���f�ku�C� �1M�_��H�䬶��;1##���/�-3�u�UP�i���JC^�����(2*�f|��F7�>��H�bFG�5P��Aol?����	E��o�,�槬��)��8����V(�J���U��I�L�0F�Ĥ�$`��3EJ��s��'L0^1mg��7#U�`lj�Y��4SW�c���W��l�[�X�l�F�ir��2�rV����!����$,���9r��%��I9c�]P�"�S�s��䢙S�/��b�r�jO�z� d�!#��Jz�����4��&�M�ڲ���B	DL�C�9��J71�^p�6 ���t�kZ%f��i � ��c{�a����Pd��d�8����h;`.�|�R�(��c�
{Y���1X~p�v��Qw����o�R�u�� @���Oq��??� �~h���[+�6�k����F2�-�<
�(���7�hp�`=;�y�h�L[A�"r��*�d'r���n�,���B'������X�-��;Vmjtc��%��4Á|�ՙ�@��Tho�~��Iݩ$�.Xg� 꾐s[&<�-�"��6
���C[�M���ƪ�?`����wV�o�-�5�W��Yr�d��
4�)��C;0s{s+'j{d���/���dy�i�
�m|����4����M�~�H���=�پ�^�I��s�!���@�N��)�t/�CD7��X>$Uśg���yv���|�3�a	,_ֱ��n��TH.F�J��]~����5�.�=��U�y	{v+&ɢ*6�����'og�z�����IO���+�Q*��qw|����+�'�B����B�$��%^���`;�Tj��c�`Ϸ�7.�Q�$�w�D��N}�XQ�� �&��]�ݲ@Wv�R���D���O��'��'�;�]7PC _��<r��ɖ)��Ud��s;)�Wn�~|��.�mt�N������);��O��c����.q�����:�oﭨ�HX�Dݮk��n�H6/�\��9�
fA ��@C%P�}sjQ��XZٗ�%,�����O7S5�a�N`�q�A�>G�CB�R���L^�듻���`�^�@1�s��4���7����I��]�g�B3��i;׿ ����(��&minF ڱ�W���R:7N ًӞ$�0v�_|�}ᢲI��u�v��f�QxU��e�"t/d,nLՏ������+`��NA�	�[�Jlc�h�%R%�0yd��S&�Rw�}~� �qh{^|\b��P�Ӱt[��P�0������E,q�䗹�Y�<�7�Oy�QƢhv�	T�"�o���s�R��	�&�t������h��`Rdq�:�
3��ʑ�/"WA����|�D��B�p�9C�0��I��~r�ׯ��Ӕ��0�=6�s�����{����[3��8�]FV\jH��
��r$��*���9�=]���YJr�~$Ѽ�Lq+�U���S[>��FNj��ԇ����8ݗ�J��mB *K�fY��G:���$�F��L�縗��R˹>�����F�������#w��n�=�͂%3��z8Hp��(�x��_T�G���}�}�Lhs���59*X6���U03o��DBka��vg)���[��~ΐs���s�US-D���Լ�'���hJI_P�k� �F.�`qwލ������Tŵ�|R��aM��I�=�5�� u�x� ��~��os��<D� [:��~� �C��[�\����ÉСI�Hw����'p�y��茦_��\Ps�XT���[�h[ܱD�B�����+���g)��>���y|g�k"AT�'��&��o��$�?�	��V�R?���AN��F�c�t8w����M_���0C�98RsXs)
L#W��c2txiG��3�4چV�W�0��pA��3�H )`�
M�����>by���]�&n���)�/���5�Bu�@�+5�s��f����NeN��+`B!o?���'�	W�$e��Y�l$��?H[�l ˈ�G1�^�e�9+�[yP��/X��cE��
?se4�� �et�q��hD��Y{��*��cZ7i�\YPN��̄*�Z'�5,�툧�I@]�x۩����Oe3i�*�����Q� 2�����9�c���X���N�KMF����&���˯����Lĝ��a�\z2���В����i�M���R<��WjT�"��(ҹ���@��Z�1	�2�5��2Ec:/��S�0�H0��$3��搩Vo*4�Om&���V�rǶv[Ƴ�s͒RK��K����4�3N�)��a-�"�M=��f�U�)�GN|�8!?��ǂx������50VX�Ay�\s�H��@�8<�i�e��p�=��� �ΨK6��ɽ��������[���L���Q��P(^�w�`����þk�����+´r����yEN�`�I�*wz\_jL��~z�G�
_�	g�I��b_kZ	�@0H�|��-�$y�h�oG�5�h��`C����JvO�C���q1Ҩ �������9c>��)0O������B�ی�<�/;�G���Z��|k����2�C��\g�o�.y�r�Ӭ3�Z".ZƳV$M�����|>%�Z>ŀV/U�p59L���U����L�f�y���h(�bb�Q4�شuT��ov�-���Ѧ�n"@����IR%E�H�| ���ay��xm�9YM�Uy��]�����c�f�&���*%�Y&��=f�����K�z�2��Ĳ�q��]���]�1
�S��Y!�Ż��O��%����Ȑ�.3r��P�6�ی?$]�k[=L�:}�T���荔���>�">U�zI��O#��$]�Z�)�% � �;�G+���p�a��������`(����Y$�;)iN�C�ꪮ4��p�w�ꂎ�y�Nя�>c���z�n��0?�g��4�u���E3e�[��m��g��r���m�dDme,� C)���̑O��^�b�gr;�a��"����V�FӋn�����T�U ;8��&�2y4�4 ^��e��,��G�a7��U�Ҁ%�̱e]mw�Y����d��ʶ�C5�����x�ԟ��Lyq`z�M'��ܥX`{��qx�^-��riH�O��ʀ>@�4�U��v���9�o5i/f|��-��0�'�E�6#��1�%�z��j���YƊÃ�X;U��)v�؞��ߑ�u�⑕28�u��>ˑ�߭�n�z���J�8n�弾�Yv_>��O*YOa�o2�'q=��*+��G���@~m�&A��`�ã7tO����t.$sɶ �J�Ǘ����G	� �����m
�bA%'��`ҍ�L�uz?�=3rclK��(����[)8f�r���qU)MCu��Ѓ��騕PQ`�;�D	�ş��S��!���L2�_��Ύ�Z-Ok[g2�sN�aά,
?@8�zI`�K��n���PQ����=�����̇�P�*_(9��۔&�� �. .��뗏!�zq`���݅&�R��3����o���������p�?�)J2r*����JR� �w�5���v�L)~<]3��I����aP�۝^C��-�7сd�P�3-�L��d?���Td���§��fhō5��H���n��k2l�-��Yj_��Ss��J��P]F߶�ǫ�	kϯO�: �Z��,����]��1lb�|Z����֊l'@oed��rm�U�A�S�au��+��5GF#{�g�z��Up�>�ͥn��t,*��[{C
3��ڠ�Xl�=�>�XEC�B��K=��A�\���F�B�Rؾ�S�1G�ή6�P�%jؗ�>U�z��!�/���'�A��(�HMtW�f�.�?�`��'��jH���2�a.z){��A���'7k��f>.�����Sxc+�꣖�d^努\���R�F��Ӵ��dL�U����	�P��'���~�"��������r1cR�v���N͉Q]ܥ�3�?|Yn[N�Sص
�A��G������7*p����Q�>|+�$q:��r.`������A2����̀r�G<�L66�E,y�.f�M&7� �=����o�+[�l_:1�;�	�%H�]�W�f������������?�P|��l����E�uu_�d�$�z,� ����y� �rY-�� ȴCü$�h/9_�w-�^�U{\t�P��p����*�o�7�<��n����I`���k!��͕��:�:E�аTs�Af��ZonoÙθ���i�о��ݣv���U�����Xk�oV{�:�Hw�꣼�Vb��uK&�Qqq
s8k����x%'d�l��;,)�����G3�E�	U^ց}�ɨ��H��D&�vm���wЇP��[h�g�{�D���t�RF(f`~<J)��E�q:i���P�	�)�_޿F�]��pր8SF���"r�|j��R�Λ���|)?�o�.)�D\�(��H�	�L.���"���f�~±"�6[zt%��Յ|)C��&g�LI���O����8ȡ͔U������1��ۇ��/����Ь��UA�)��,��B�O_���z�H��k1^�Ɔ~�*[��Ae�ΈO�o���}V��Kp�_�e?.j�N��gy?ӧ�2i�eV0_RvB˵���ї��\���� ?NKa�D,=C�
`������Ӂ܍T릸��������� C�t�A�/q'��r�9�1!GP_.��0�&z�������:�|�1�Ty�a}Yq�sƅ�L��iǌ������.����J��Y�K��,F�����.�x7��l�#6+T
ੴ�	S�~�s���2�	o�AR���L��<�|�:�I��N8#��S��r�@b["�%�Z!��=F�8f�CF_3#1��y^�w�ڭ���ޛEw�TcZ� z��P�А<L�m�$FM�̸CH�Ŷ��;v*Mɻh-^��$>>�,e��;$.�Ɓ�mIv��P:4���v*w��~{�v��6c��ןvfn��JV�^�\WnӿP/ؘ�#�pqݝa	mϖ]n��-�ƺ@b$���C�	��ֺ�Qy疩Z<��9�`K�b\މ��J�x{j�б��j���5h(q�uH+����2+8ц� ��p�1��N���� u���7�'����*^7c��nbg}���D�m�Ŵ��h<G�/(��I��*{
��YG� (`N���Ր^�lń���hi�ݞ�܇�mt�]D�r:�AП���TT��h��/�B��/#I��Q��Y��,�;��������j6������0�yU ��U���h 'ͮ��o��p�p�g�ovг����������6�)��.ϝ,�x{߿,��]����#���m�y�q�<��O��w�����5�i�{��y�t���.=����_x�����j|]�\������t�Dv=p�%��5t���on:P���o�㾸\�3[�:�����,{>=���H+� ��D�ıvP`B0 l��XI�V�
�Pu��=x���N�܌?ly����������<O��~ S�͸�ӂ�����S�\�|+��Z9�ѱPWx#����Z��!�� �������BT���I��_K��Y��M�.]�p�����3�\jAKr��c.p��V��Jg��%�����U<��7a��^G:�T�3�FU�Q���*}�^ �;��\C�m�r��`�F�<��R�Il<h� �W�Q�JT�cD2\��TS8Є�W��%���z]R��N�߭�o+��FT�ZZ�v��y���5ņ}�	��n&n�T�oN�!�1iø���<f��j���rP�n���C�1�0�jS2%�n�>{7�k�4Qh~���[���W��@�Q��h�)����������`>��;1�J�>VϳVV�m�IÔ�e�I�>o&٧1J����V
�vND}��Պ��A�/��2A�T� Q�0�:x�5�Ob��e碠m����B}�h�|�`���bp�P/�*�����WO�!u4�^[b:S�t�v����1��Ԕj� �N�א��wN��4!��\ ;�^q�B��`���h ;a��ʞ�U���ޑ��ílY�9����C�!�5��0"l�:�
��H�3I�%\HI�Z\���R]�¼z���D%�"&�k똩��
l����6���p/��������T��@��}�pnG*���6�������n!��J���X�E��r��nd��N�7��i��Fg�����hZ�'�U��"(}�~Xv*�<w�h^�!zN*�恊�%�!��D��`������u�)��lct��u��~�8�l�6����p(�k��A���2��)�v�������D�`VU�#Ah��u��g�lQ�<����	��G sׯ](�&�'0��$v}�y	qA1et�����SN���ma=��>���<������#pZ������Q��`B�ە�-�ÚWk��$+�ԗ����*VWM��^����c�}�} ����8_�.>B.!�ti&\�6����,󺙏�$}t� =�9��������k,�OYK�ڍ&�n�ul�ˇ�\��-�C���18&;�v#<���Z=zXV���*��?��E�`�N�p��$S�XgpW}����Y6,���W�xp��x)�	i�HVtYX)a.����n�T=G�� �0J�9�e�k�j8Aɒ����:�@.y�����t�en����D'��C�� p�����8"vԹ-0�`JT�.�:}Ƨ0���J#*��6��9F�V�� 89B��K_��N#�}R;���N��=��c0�6
�����1;"#��}wF,�:�[�h#�qC�hNX�������!��e�{��	�8!ccy�۔��뮽�+�obl>�`���3%�j
:@�2C�f���p� ����Z����r���EHq�l /OԮ��eF�پ��<}2b�oM�
\�Bt�,�>��q���U�7ļ�yg�v�O�,���$^Po��ݱOR��6h��Rߑ�����1�}
U�<��t?d��R�|�W*\�p7��q5�[����x`k��^Ǚ�oXT��]9�/fq=1�̩o��M�ɜ�,@�I��%2j���*�c�:\�?�9�N�sY�߭���XP�6rd� f�����6��I��t��F�_�jY��? q����օ|�#ʭ#��W_$Cl�U�ަO�����b�T�p� �c�*����[<�4�xU��a�`o��}�����xC�3�\:�H��E<1��L�,@!u��g�2��͝6�ܮx�{#cz�3��n�^�U��'59)!�-�3~��s�$�C�]���@hgm`�>�'Q�Yn���8�%'ϳ�>y��v=a�L�8]Xn��&��Py
eZGK��q%�P��Z�yƸy<��|@�ǒH�M�RFRHt��F���J���k�/D�{xe9���>	���j�*��R	�6�h��<)8�`ā��lإd�7�H��H���>.��;+�*X;M��؎7x�h�R���v�!t�d���em�rL&>��:m
P�콑l�1�z��q(tt�xq�G�wN���<�/�wթ�T(ւ�Cr|��9�@dH�54,����͈Y=0���(�0""�p���di���9E�1G���`۰;k;^!h`K޽J��zٲD�<Njs��6d�����1�$l��U��V�JYO�^�g��l�g�g[\�zW�9�j��f��9RRL�D|Y�������&�9�k�����&�v�C�k����� �Jh�h�8᣼v�&��A9g�\<���r�_o�+mĳO��n�T��dOe������I<g���D�Pw�?������p��R��Ώ_�E�B2���6�O���7EW;S���Ҿs\5�����)�I��O�>(�*��=�_�u����V���'-E;1*h�Ife�l��g��;����B�0�'���9B�X��ۑ0�勞�)�0޿|{P��(�m�"1��� /�Y��
����I\.����$#�ʈ��#�|����}'}�0�������_bʳ�h�Ӎ煖"Q��#B��)?����Bq��3M	�rT��?P�P�߼M��rү@�GN���މ	�l������ƁV�=@�ϻM�J��9^��.���*#���6�~@��J-���Q�P��y�H��<��8�Q2�ˆ�n�=v�E��dL�''�&�}͘p's�ەhǳ���h9gm9��(v	Ӷv�d�s��mx�.��;w�=��x��pƒI���6B�pA>�B4���j3�o��?�O��]��D�{�<�4W��ߕ9�m�7�������Yu� *�4��g�Oʫ�$Ék�L]�d6i��n|�v(r@�,��#�FX;vFq\z:�Ql=&���1iD�:.�a�D����/X�~U>��'��U���E�hP0�����B7��Guk�>:��N��fD��z&:��8CY�%���-sߌ�j�Nc�!��H@��l�=�^����må���-�P9
�ù����3h��jTBĕ��Ɖ�&jA1�҇�[�9ǫ<�:� �G3�4�c[�2�y��8��^�]��҆��X�xT��)�����k��{��H��r�7gm&1}��	�g*�fNI|oIzP�穣�i��.�`��D�nz�\�vZ�G��#)�rvJV���Qy6	��E7�m��I;��X#�dؘ�ͧ��3cy��2���Ds,b������mMvq��p���~�����J۵o6�SgD?i��`v��`l�=ނ��5���ƹg�~��z=��gcu�Zy�)��X^}�jͣ !3\��f),���M��Qłk�Ŭ�g��.#��۔���	l�?]d��a`5�}?��<��l4L�\;z�u!�������g�q`*��hm�!�?�N�LQA�\&<E|"^�T$@7�t��H�tN�w�L&��@.ؐx%+����}$��:e��=M�!J���6T}]�rg��n�fn�����M�%w5!�3�g-��y���8�^mA;��Q=P��T�����
Q	c�*�/�9y��$/[jt��p�G���p�놡��L:e&��V�n�U#�¬���K�����4�^��I�η�ԑ��(�Wҏi��9K�1���f��W(w/�Al��1�{�#��~�%ɺ�Bܮz�Tڲ�!����Er#X�}����ٗ>X̨pe�	������Ŕx�HKP|/�`��������zu�Hj�s�)=���ˎ��LB}R���V��~^|4O۪��QL���h}�榅Y�-�v��Re� ���:~�e�H�K��Zg�T��6��A�D?����eDa�&0�QT��R����L��	y�ǭN�pOtu9� �uv��O�N���~Rm�<h��T �0�+}������	�X���{Y�����|u�?sѪ���ʇ-�dd+C���u� &�k�^�2��d�*%-�>щ8�;��]�1yS�ݧE���R���� ��&� 6���>����������C]۽m\+% c��B02��8���P'�
7|{E�M���|�ğ�3���u��"���ț b8�����R�+F��Y ���.��vCƣ������E-Y&�I\g���$�#]��'��c�bb��}$��	��A���U�mN�&���	�a��E|�z�u��&x��KX�����E��s���#s�ݎ�9�ے�������^�<�s+�-
��U���w�{�!ĝ)���颂[��sS4!�=�{G�{�V�U:z�W�V���BB��a(T�(g�@O�.�m�&�0=]��j��ĊX*���s5HD�= '�x�K-�p�<{:d���|	M�o/z������ m�,��3��K�n�|A�[������`of�d[�*7�x�?BQ2� �sV�r�X�}�;��n�C,ķ�v� 	�G�@�t~�B��z��� �<"ۜΟIv�'@ͩ=ٱ5�Ʀ>�8p9��U���70��(e6И$'��Y�t�D0�<�u�T�Sx���$�+���g	"
^���фiɃ�C�#r�L&�xm��>f���/a�+��t��O�
�����
T�?�5�����C���;�?������ԢMC���C���a���E��d3Ʉ�M PN9��P�1�m"��倽`~�p�5���D�GV}/cI����#�A(�	���K3'����N��l�TGK;A��2��>��q4X:hH����5��j)@�dyVـ�y2�>,Tv��/���6�1EY�`�V�A,���/t��[�^]�V]�z�h�%jbHL:�Rj�LoɋES���OY0�Ѯ@(�R2���$�_��h�&b�������Ȟ|bШ�DA��S�v�0z��o��`���=g�k��n�!_��>wP�jq��<q��g��z�X�}s�6�z�B����Db]����;����ͥ����g�}2�:��طc|A�\�J"�*���
LIl�m�^T��m>�����Og��3X���s�L�
y����%-t��A-��BHfb^�m�Ҕ�M�˃U>!��!���3:N������#����A;��ok�9ގ;5\`�J�ZW"C�֊�o����q��ْ�5�*�:ɂ����סC���Y���Ry�=��'r���]�C�}3�I����ʟ!$���#h�Y�\ȩ.k�V�"+(����E�+e�V�˗�=vTq�������.�Z3�
:�P�G����h��)U��!�E4q<�77�XO��Z#�����ҫ����B��d��`�
x�I2���׭���0�g�Nzi�䲳Ǘ�"!��U����ɘ���U��`�k�O+�gӀ_"����Ҋ8a:)�d�aB��mU�ylFv�>��x��?�,,V�8����,A�=|��}�����f��v����%AU�& ��"�1��|�s�<�%��*j����f�:{��9�CF �u{W0��t�S\���h.x�,\���O}[�c�x��ad����x�M�s�����YU�13�%��|� {9�0��Y�
МH��]��,��4��І2`��a��M��������Uj��d�\��5��v�K������w��LUs���!�K��b-�q>6�c����9T6����e�Ock�DwR�K�Z�p���!Յ|�}�� ���hd��G�@��:<�F��k��h�L�Z�+��,�r�e\mJ� 2�U)�F.=�T����	�	KkH�SST@]��\g�K*
Y�^~���Oz���
���	d��Y��G�'�"�.�������[��+���M��gv��Ջ�Ɨ��9M&E�)�I�W�m��Ӗ�И.�>I��a@�c��}����qK<vl�tt�{�R0d�جZ<���B�� �J��Q���|�C9�u(����2�k��X��^�/PZ�0�����>M����o�OR�F�Oz��څn '��f!:a��c1�C��8��r>>=��mq�QqGdj8���&�J�����-E׊sLJ�KA�cW*�;+2���;p}B�{�����T~-��S�cu�������Dh��?/7��|y���^�9�A#��~�f���?N]�F���ߥ����w��HIU���@zB�)RE,����=�f+ił9�i�@l;���h%�����"�*�mʽ��o�CCAՙT��h-�h��}I�:j��㊑�4��[���@�y^�̿���6у,�*qL�������͈=C��F����u���C�q�.�\p��A*|���U��IYXm�p�:�C7�O˷No喪?�2b���/E�A�
�u�y����w�A|�|��E���l}��7��Y��VŜ�W����>H(�!_m���	E
ĭka�e�t�����s���ji/ '�p�RT/o`�	��q���d�J�DnR��%u��ڎ��
Ƃ��f&�zU�T��ɕU�9�Q}LM1�.ެ�J�k�t!)�SG$
�J�J��9N�)Gx�7�����%��Hy��z#��)�1c7l(=�C�"�$A}"gO#���*��$��Q�kM����75�M����.@�z��*�U���ԯ���}s�*�@�U?�'B#�2�����g0�8Xl���(���frF���
��&��a����fX-�Y���Bw��c��.��Yi��7�v@�d��޸�(eqep�Ʀ���l���k��L�)1wB"2�ܤ3^�V���k��
N�Aޱݎ�f�"'���B�������$��U[6�&�M^~��P��C��^���l�/0�U�AX�>�C�_��Εd\̖(:f-L�+_ظ!%��9]ɳ�@uW�mf�23�ުƊ�y�3w�|��%]�o_}$��;�t��V��ͮ�5��L��?D����7(���:�����5O )8�ԧ��0H��a�@��\I���A����ҵ����k��xws�O1�#\*�۪�ҹ�=���XO����ZC�ƞ� Us�Z, ����� -�}��j��:%�&�]!����P]�;�V�Z�ء�FǓ�.$R�D�(^iZq�L�Z��k%"C�f3���۪��9�����G��h(6�d�7�\7�ܟ��Q�1v�"�bX\@�\��-<x��Y���x�9��l�!`c�7ʾ	G�F)��:io�Kb�1��<$���q�ኚ��[z7�J���5R-�e!����%NB[u6Lȁ��cWP���M&�����V�]���b^��t�œB���|٥�b���&�рh�53��K$Mv?)&��x�V>��U&@�8����������YI?<��d� N�J�z�u���h� �'Xխ��4iwe�j�h�MX􆗷Z}�.ұ�Z��.�G��{���B<L8��EFj�S�:d��* +�5���/�XH�$�s�9Y�J2r����#���/���f��;�`�$v��p�<��W-���}�lG�����83ߘ��j^	F<����;MeX�n(o���\�|L�{���dp�2�]+O�fm�u��C|�%�fS�o$�:����6
c�����ަ���'父3�e��0�q	����ǚL.�J��E\��x�]Βj^�a!�O���"D��W�/8��?<x� 6W1n�I��&�X8u�g��z�O�}p
�����e\�"�}* :���{���j�`��� ݶs�ɪ�MN#Aci�e^@�'����'N=2�����Pw�Wx42]��(9G���ߞ�<�r�gGT�3M��y�����R
�T��d��Y~�Y�:�V| ��$`���9�UN��Q�\m�Fg� ��/N���I;������y$>�Bl� p:,��Zɱ �����dS{�3��kj�h�?�-!jh���*�'����*��)n��o�n�[e�t~5KV�#�̎[A6�J#��F��8��Yoo�>�l�I<�
��/�l�ɋ� m�;�]h��50#�rq��Q|N�]�d����d��2���]Y���D\��@��g@��U�� .͞�D"*��ʴ�D��C]�DJȬ�tm��ѡ����K2L�u��s�R�L��]�2��k8�Ш*��C�T9�R��'[��9ϧ�s���ۨ���M���V�r�J�Ʋ'2��yyl�m�����F��7��a����02���{�W�^�t�O<���hڿ�Z���_��	���ܲ����\]�Als}���軀8�0[�����n?]!�e�5w�ˮ������B`蹹���!��>Q'W�䫮�o$ܤ�Ҟ��rgR,�z-�5����=&�
1�/��3��L���Aw�g��#�J��2�A���
�p����|+�&���T�^LnK>�T��_;%�� ��p��6�\��o��-J�'n��,�)9U�3�	�a�O;�Cz��9�����ƙ��2�{�1�V"XL�HN���=�u-K�0\<��&�=g���ԁUc��C��V�1����fi�����Ȳ�8ݯ^v{�fz��lX�%jpʂ���q�e��t��B��?�a��	���R�>
F�i��v߅�<�Y2+#^b?�9�+l7�z�8G}�%���f��=����S�&�{��P|�TNv�.��y���\���A��t[�rv���P�+	~��e�J�g΀�V-[����8]Q!,e�I�L۾��TA�xɿ�I'WP_�6�M��MWA�k�x��$��d�7��s4��OVx�}��!��U��JO�Ũ=�F������H�2
�nC�xn��1�_��+Z��=�>�7`���c8�簽���4��DGa�u���qe8A�f�6�`��_�n�e��X��)��W��4SYEPW��ȎT뀭�7�@b�(H<
��a�oA���ų��Z
�'�U�d�~��$�:��VMu����Yq�
�K�$>����!��Uv<�>�����3�Ko��"O^�$ZN	h���U��@���W���Mr+�kSyk��?�uS����܋���ߟ�9�_!��u��E�֯��py�@��yvp�y{/j������o���X�݃�
xt��AB���n��!�A8�[��z�ҵ�.��7r���,��F�I2OǣPK��{ �f��L�����9>��bd�$}E��?��Q���i�Sn}c)�������HZ�sz�PRU�P2�ߡ�������p+������?}x�5$���i]���wA�e�N��V��Vd��*C�7��z�#ՑHC��!�YV#�����:�SV�2����p�f}Mj7���%��)Ϣelo"Z�4猚����PZsT.|*j � 9D�rk,�?V�� ��#4/�X)�ރ�L�O�G+��ݾs�T�Q��J���x��`!�R�
�}���i��X�'	��}���b��Tl�9�=�d���#����N�)>Z�9�{�z�?����5���2ʷ���xI�oZ6k��{�2��ܸ\�瘩�����f��ƹɵuR��Nuh�]M� ρ�g\�$���S�?_nt�Ƽ���y����Ab��4�������s�ЋK�X�ev�D��4;��I1��Uz�~� /,Bq�t��}�{�����z�C�5HĪ��oI�Y(�#��ukI/�lX /�7��+k Iv�}1,�u�Y�jZ�գ�n�w_@������fJ�=W�0rYdF���|�`=?���e��( ������(��=� c	xˇKl^�?"���7dO�@O��j�8 P7Y��7H˓ ��x��R#��I�C��� �Ɛ�w��~[<��!��;K8Lv+������|���]KD��Z����]��#`���X#G�0�Ʀ��î������r_���11ĘI��|n��/_���y�#.�L�R��=�r�GVVvWL^]��U}����p���@�}��l\괂,����8揂�%�bG}䰇e"��/CV��D�z��߻�斕5[52�y�*��1�a����O3*�;b]���
R�N8���
�X���E�|��f�+�W��r䗹PW� '}'1},GW���Ek��,�'�������D�X	7N)0�$4ۋ�3����M�����{�_��:�	���ӟ��_^|e?��6J�b!,��ɋ��,S-��i���\�W���;�N��xP;�h�+~�����{�$,��-��'��:b&�i��O6T�x�ZHJEd7ъ�{L����\m��8˃afiV��
 �D���[�>֣oi�NNa�V������<�\��J/X2!��O~���0S�����33BL��km�?�;��
�~,b�jA6��
w��\�6��d����O�ē���ո��n�cy�m��X&��q�p�bz�G�}v��r+�$�џ� ��QA��J�D�Ntt�[�s�⠄^@;~�'� Z��g�ҷ��7�)�sFG��	��������s�hQM���R�i��7���B�iaL�e�t%���>����42�i��W���B.�O61�K�ĳf{V�A���P�2���`zm&�s^dîK`�֦ކ�	`e�Jd��5�[C@d��C$���E��»Ŏ����q�j�YD����s�>��z�vN4����-Sw?��F������нں��34�.��a����������[6��q�&��4�
��
�ﭽ�6�R��5�����}�c�������5S8`�z�R�@�R���9U���#w�ѣ�y��@��X�_�T���HAg_[���_��7P!�y�?� �տw�����ܹ�.Y��."��@'.`fh���E�,�&V�h dg4X�ڢ��G����mv�p���!;���L�*)a�Xo�1���1{�oX��z?��I�c�����`��KPs�bY[�6z����_Q6#�q����)㈁	V5[��=��ek�4Q��SZ�s�-�j�d�=��gb�E���槦��<�*��-��r"� ���i*���%�;#�0��dF�Z�������A�N�#�=n]�ʲ��k	�9�����X����$���:�=��rz��+������mxӁC�ݫ0@� w&�yڅ^�&��h�ڬ?m���P�،.Q�	�������_S��|FdKaY���]���o����s���!�Н �dEz�g���o�5��|���M{�_�%F�#M;PD�+ZU#��O诧��gEmy�Jz�kWS_9:Ʒn����ǯ|��@��}�U�E�u�*��bd�%C��[�-єPj�K�`qf@Ư=�6{L�Ȧ�-�y�d��D��;��V���斌t�A��8]��oɽ����Dv������"U�{�������,�G�7�@��B�ՙ���zRݘ��,�������>��~%Z�xS;�ִ� ��E������ܽ��y�*Y�}2d�GuՀ@[��BA�>�� =]<��#��p�&����=������Rw�v�_ې(M�
���|"Db,P���ח8�� V��?�t�+�!�f�(>i][�I�i1/�h�3
� qa>�A��{eM|J}S*?�L��?��0��okpD�!�p2���v������j�_�j2'/@|\�����ڶ�����#�t�RYm�6�fse�{W�6>%�]o`Uz�vo����b�4��X�����l�F�u [���$f�+����;?��BO�ې����7ogO~�׉#�a��M�'ń,4�S�G6��������� ��L��� ������ذ�/��%��;��H�ϼ����D��_^Cx����S���K�������bJ�9�*~E��L�g�E_ǟq�ؠ:��e���x�v�;V�,�a/-�D��}��A��2���T��1�}�T.k13�ѨN*p���Gv��p-�b�{�EK�B����O(]��?L�q���؂$��3$Yh?��ۆ[�h��Z�=ð�m��*�fl���ZZ�?acz�싽�S:�����yVkG-C���ڦ]�8�7��js�N$yĢQbẛ�u8a��ZvsjB�A�v�-�F�D"��4_�1#���\ȸ����hL�H_���kW0Sy�K�x+5���׉����s��s�~k����8t��4u�V��q\�~�^��g�P\��U����Qw�g�����{����~�mo�����5+H=`1k�2�H������c��U� ��_8��4�^�<�@���l��:�-F]@�&��h1\� 6cl��8O<k�"���0!bz�D7:w�$�M�4\3�l�<'� h�N��#OV�aj�����v���֗-|`�D;��S���eb�%Z	#"����=j���P��%_�z�X~fl_��i����F�p�x�o'g��01�m4V���&���)��(O�����5���I��&���80�}J�w���&��ޝ? bc�|.�ߴC#��}�Nl����d{U�֖& %�G�j��B
��j��[�4�����Ka/��r(w2�t~6�.��u�Y8�*yw\��w<��T�|�����VW��P��� r�|`�����'gp,Q ����j�lT�b���I��g��Q9��1
ϚS)s*���F�N�ߡ���X,*s��!!b����MG��ui�h��jp���_ZT'�/�榸������m��`h��� )�|Z�����41ہ�#�N�ڕɣڭ��z�jF��w\z&~��"�R|��t7M����z�Ll�V�E����L�$6�N�v�'saظ]�q���զAy��1ݡn�&�7<A�z��A;�+Y��~�[F�$g;
=�%�e�ooCfŚ���J�ȷ&���\٫�6m{^��H�d� ͓�,���s�Wu�⚥!�@�Gj@���O<�c���� 6wD��A@�9�s�F�bH�?�?������esYZ����dV�}% �@�Sig�U���Y��2̭���^��0�ĭ�@����*W!� �oZF��n*�X�b��^��x ��<K�����������_���0C�Y�GC��4�K�K�&�*�C8T�I5�Y Z!SR�5�}Q��[�LUŪn���7!ժ �ws�t��#I�ě���I�d��r��v�C�Wu�TYC��N��!,��(%`G�9��z��o����4��R�%����]X�E��Jو*�\�3�٧i�6�&.q�f�" ��z�P�A�tZn�������
�f�0��N�"����J�h�%9����/
j	V�\u�R�P��
W��i^��G�s#���Xȩ<0�l��q���$��|����R�}�˴W%K\4kǊ��M# ��\�O�@2@W���hَ�!vQ��R\\�@Τ� �[ަӤ&\�O|37/�`�z���)�nr��D_���lR�cy=���
�Q'<��'%��m�l�S7~yњ ���O9�4�G�FjQϵ�B�Lq��Sߐ�x�ZV�uܱ֧�H�:=�;����62�Ƿ�F��@Rd��LT���Bkg���v��#B�ǋ^��ɴ�i��bj��7|�wd�]�}�Aʠ�О�� ��𛑍&��f�ܓ�����4ܷ�
��RE�Ww�x�ɶV���������}�=W%�xFw��\`�)!9���`���ı�.(���|�-VD_+g^r_~-;�&ȣ���Yո햒�Ň;ܺ���ڶ����J�9a9�;ih?�@��ѥP�! 8�D�r�~�w6f馷6��9�.��kg�����rmo�O
;�BE-����d��3g���I�xX����R��w���T����2
���_��fB�V;D�5����l�B�b`���v�ua��'�;��
v���`�S��:F�
��b��,�r�Fx����R��� �i��C��;[�AT��s�'�%<����q��v�n?�̥���;�W�S���}��/Y�w��*-kL;�-/�c�;0�c��7��?TƺkcJ���&��BE�7F�25��]�v_N�;����Nu�r���/)��	qߞ\ڿ,}l�nmլ �݄���ԌR�n?CUmx�������Ge�;��z��rC�Ge��8Fm�&�i[�w�eeU��PU'
�Rw���FA>(^$bq��񼰻\4��u�_�9���I)h@,*�k'����WL{����`�4ڪ�2d�n�l��{jG�Z�7K>#Y�#�R�0u&�ﷃ��_�����JI>��A������ne�',3�K_��������Փ�AΌ���?�T���r��+)����b��	S�4�\,����K�Ko����{ނ-`��K[*X�-������od��� ,d�|�Y��V�Շ�e��Xj���6�wD��/*�]��Zݎ����*Qf�j�-���L��K@U!��sӑ�آ��CƗ�G��
ѩ�@����2�j}!Z{hDfL\,���t����)�=�'՛G�
�Sպ�?4���ʐ��	���}��ͻ��*�~�)]�n|��hHޣ:��#�T�v�z��+��DQ�c�
����r���vܽ���xa��eh��l��!�7�잞��M�K�{&ʋq�$=Sb˼�ξ 4������I�}���7��4�����_���c�ۢ2�A���<��Jg�1�g���1�C�R��.���.m3F���k0�ؑy�V�M6�<��qT�U:�;�ڂ�3x�X�}��� �
W�)E���OWA>(��~�������I���0f](��6J�h�*+���'�]�0VI�g��J��d���/���9A� A���*��s�KG^��f�Q� <�Hsԭ`�� %��g�ja��,)�u�#�HR��y.���<>�+1�({|�A�խy�f�D�ּ/3L�=���:EGL�9�Ѷ�ec+ ���%�@`���j22���y�k�����wO[:[�|�S�r������:�i701�6�]j�qS_�&<R5X��g�o�
Oy��:O]?-Q����	��m'�B��p�e3�Qb1�Ac K��kX��)<�D|ml�1^*W�Fqh����b���Đ�K`(��L��R��DIz;�L���ٛ�fV	��c%@	X�����WL1����y�<*��
�p7N3a
o2Fu�O�/���Fȼ�Ť�r��t^�>;W��r�J�Ny.r_���l AC��x�/��uB���;٠��]�a�u�kJ����{��f��N\�b��a��x#Y�w(�MT�'s��h��"�$@l�n3��`�r؅�[���Y���[{M�%��u	aK�.��>�rN�:�o%��!�lN����ǘi�m�����ֿ��#yPQ.��_Y�5 ~K�0X �Q�����ZM�+���U1X)������j�F
f�J�Hg����l��;g�;����L,;(�0C�?�p[8�Y2R���%����xm�$�!&�ׯ OU�H��y���/�v��q8а��Z�vs"Uo��/�ms��.y���0�U����:J����^�(���C��n����hj�Z�m��R��!�6O�� ߵ"��su����dMЭ���Yg��o� M�p�5�]�2�����^���\��������֪!���*J'��V3�1mR���ؑ�/��oE	ˤx�A �l�:��sr�&�{���_eb�`/�\��\���"�����F�I7�ZdrR|�ߝ��ʆ�ކ@�;W�]��(W��0W]A�����&M���������)���rM������ko��hY�"7*���1��xT
��(Y�w9O  '�Eq&���Md��O��GI��F�J##p��u �y8
���%�t�>��ҫP��<_�{��E�F��b��[S��{�XM�^[ě@ê�S�;�q<-�?3�ˣ��0.سV��uD֫8���v���E#M���^;��ʕ�=��O �T��	Lv��t�~��뎾�{��*ם	��%֔2�	+R�9? ��SJ�e�G$me=�#�/��Ù�9cH���n"q�%�q3���y���r��	��t�D���t���\������ ���3�b���b�l?5�����+`M
i��J��(�z�`x��kf^���3��A��R�&\Ѓ^��L���AsK�mV󫤏,�,�����0�T�ߪ����مq�nDM�a���ݽ}��z���@�K�7��q~�c�W� �bGܸ��E�ӛE4��4��s�f�����Ì�X�۫(cag�}��9j|��;U�V�~O�I�܍��Q�X� ��&��yv-ƛ�o*�������4�˫z'L��Lm�S�OJ�.7oV��kHB����u�r�>���C��K��U)Q�~ͭ��FO\
c��gP��0�zf1�AS ����愩@�/�4��j�(���3��|>��!VK���f�IxƷh�B�b�@�O0�'�c߹�|�px�����xħ5��9�t)�Ju�D�R3�S����!��C�o�'OReZ@WX�'��wL�c^���]��ķl��K�ܻ&"���}HRO�?���63���H�t���b�iff���Z�ݳ�Ua�<�e+bx�%�ϮE�����tZ-DR��D�~ĕ:p{?)��i�'���V�mL��wѭ�#h��=�N8 #BׇI��ݡ��ɹ�{���M�ǩ�{[���vxJ��dx�}f6���4��1�aB� ,,��
��0�Y=�*i��T�x5��h�o�e6]F�]_�t��"T
}9>$�	>��y��%�*�f�3��K��������{_u�������~�a��eςS�j��XS���[o�Ud�"+��n�� �+���'e���P�f��{K&��`��cv����x~�	E��v�6��x�P�����Ý ���?KM�����Ue�
:I�G�b�8�}aмs�D}?t������4r�jؠ^/zaU��x�����븘r���pY���SiL�	�ha�&�t������漐� )p��®�(lo��Ae?��]��Jdؼgr�q15�p�h�߅�$�n��Ҍ�8�!!�C�oc�����4%7��(�gY�� � �6S� *�NP]\sT�+�q��<%Y�UϦ���K��L��g>j��c�>P�9#̻I��umr����f,��E���._��L�F2.8�/�Z<����@e1�ȏY����Xq����7��%F�����rvt�Ð��'4%g3�W���H����4A��aRyDP���}�[:�3�zԚ�V8��Q�l�ԋ�����H ïg9B�z����Cck˻q�lSf���q�ڜ�}���t	�/��U6W����oI��}WlN��M m����p�O����z��:��u���"���I�{i��XI�3���������������(��1=��yzw�*�g`��@�B�V���:�ԧ�W��D9���)��0�gvK}���~(�l�?(�7��c
	��z _wVj�%րaո�I�s����я��`�0ĉ|�q�:KL��2ch�B���X�{��J&�S��X�j�Ko��J���ƀr�0�Q�l��)z��R2��_Vu�ec�g�|�l�g3�u�|��w���p\���A����p����
���ߧ��2=�x\���㞱9�D�v����pb���z���/lwYM*��/�Mnf&Z�?_O�k��`{�����{BX������ވg���9�O�|;R����xz�w��e������Ñ��ޜE����|���C
��)�o�\ಀw࿧�x�
Y;����ƙ�����e�34&8�^QN30Z)<�s�������c�6�m���f	���	�o��h�=�h��H��[�G��>�Ks��=��W�}~�Š�X�¯�3�\n��b�M����ح�/	9�h'J(o�_EВz����r���r�1�d�����Z�Z��-^��5�s��>�G�u�\Pj?]\��AL�u4�m91��[�O|:���$�1B��Y�Xԉ�.~���%B�|�$�9��6C@Z,�e�����  ��9�"?��4ڴ.Y��n�>�o1F�9������?�~u�G�eܺ�f�4^��;����f�f�e�V��8�V��БN��r��J��Y���T������P��D_��an���N�Y���ψ�M8"4�)�K���u(��gżE�{�@/���P�X\�����)���Ϝ*��Z�J����I� t>���u+=�o8!U؞�ܙ���^� �n5\F�v��z��5Z�������4&I�!��7͕�%�b���<�S�֞Bp���ꥤ&�a@Ҫ˭�z��o��$3��r��.I{1&�Y[Y(3��V����w���z�+��V���q��dTu���o���"is�!���h@a��m�J�B4�Zh��h׮wuw��!\�å�ݞx��(�j��,�u��\?-��q���b#����Y��?D��蹐��`���Qàq�MX�7��[J� `1'��#\�j�!)����8�5i�c�6�r.k#��+��'L�g��B���>�E��Zi.<=�{��mƇ#�DN�Y��WeFa��n�7�ua�m ����i���H�X�şF�!JMv�g)kͤ�C!t$-}�T�_�zÖYt*�>�W���ħ<]�܀8*�݅�f,�#{��'�e&g,`:�'	a:�8]���v�@�9#��(/�_�9�����ݝ��˼h/m��-ۡ�5��5�}���i�8�W'/�-����(�� ����yћ{So$��/ʁ����2��b��v1O�|#�X�� �e�<��$��ݴT����H�V�X0X���`bD���&� W(h�p�(�3� �C�ހC.��o���%��H�~�H?���
�����17U{�2��%��]fK�M�_�|����Ga\��a��m��6$�K�%�M�k+$����9�@������x�rWW"�o�5A;K��<3���������p`Mck��m���d�1[�d�Εw�4�[;+�/�؅��:�Y/,����PL��%�8�莌Иp�4:5��ȴ޾_� s����^b5�zeF)[2B��{[8��`V�OH4�o��,�6�K�h6����� �
s�#�F�$��Z��k~Ryլ��C֪.�6۫F��U?4��Sġ�I|w�e� %��������pr�� ������`���$�K�H���\�xD9\��y�4^�e�! �~j������RE�i�H����;Vh��[�pQ}ф��'�-��T�`��OF�)iGBFp���TY,��.����#߇��!��,"X��}bƂ�G@�줆��ͩ]�	�К8v�X����v��8P�29�氬�չ����U��1�s�_�תxq?AMy�쇟"&e7X��v<�E����L���tI��C�[��#��B�����M���u�,��p�����u��{҅������X��!7�D=�w����*�3��S��d'�,C��~ޜ=	�xO�U�cu���%�w���E�M�g�+s�B����q��\3�N�u�[�b����a��ă�26���B���cD,�'!¸���������C����e2��]rPo1�*�ݣat�=m�C��E5�-z�� 1�2�J��b���ol�t�Pp�҉�@g�-6Gq*���!�sk��4G,ȏ�k�%">3�e�|����fsll���o�3�vM���a�C0ۙ���y2�	��9�2��P\sj���