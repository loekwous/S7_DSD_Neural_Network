��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`wk�~F��)١{���K�.Kp(����r8��y���գE�zןΩj�-W��f7m��q�3��=��#i������*��'����|�@���C����r�ї sK�����I���Z���?��Ғ���&����� I��L�$4*$M�R<A�ӌ���6�0��a?�w���1�s�
˶��߸wd�«]@1o�H�21�5+�v�FT5{i�2jCI���.*��Gne�0NQLҸ�M�w8�.{C�U����{�Nf�T��$SO$���p�W4Rw�F�aalZ���j��3ݸt�b%y噶i�SqC�iB�KB,���*�9���25%�-,�&�f�ʟ}�1�ۮs��{��(�0u�a�em.[5e*���C�2��Z��EP�	[7�P�BX=��o���~�n?i�퐎՜6���"�!��I��G�8l������0OH���k~`���`tQ��x��\	%q�!&a�8���ȷZӋ�8B��:��_X��5�̺ܰY�/q0��3�=� �����h+�	���&�ܴ�~Л̈́G��	Yuk0,�iM��9:����%o���=o��s�C���N?%~t袩��i^z3٭bX�>�=��{������_�*�U���SK��a+m^��S�tcc[0���tH��\3�h[��A�j����Dj#�;�f^	s+x����B�b�t?���=~����?�G��*�W��Q���(KQ�lDlM��o�#���m�>���.(;��>����b��h� �`_#}i{�!�Ԁk����%w�����E�R3�@Sx,��l��^���3Ʀ�Y�5�thǻ�2��HZtx���[�X��MDF����ui%,*Sh�X)�L��e�MA���K�fn����?.��U�U�\I ���]Dhd���4G�%���ϡ�#́X�ÁU�<�����,������[!������">��b�#̩�p�w���p��u�ݲ�4��>�$�8�� ���8��~�ҝ��om6��b���Pl�8!s�c�^�WfHm&}!'�S���hXL�^uf)@��n^�u9����z�4�pn;c�a�~�>����N�������=��r�WE�{?,2�\�ˣ3���mP�4�O+�Z3U�N�{k�x�����;T9���fҿ9�{�ѮO�z�hk#$3,��OP�����QbD���zⷈ]j�o���d��I:30�;���JKh���S�2Kv����Fh�����=V�D�Ce���$�.��QقK/h\h~es|�&&�+��~��zK�=���Z�M�˧z�.��&�:�}�[z
��/��B�O)D0���\���s�#q��R�����Q�ڜ��|��e
5�0���x���V���&�:K
(x��
l�w���).��Bn\���P��mju����vwo�ǩ�l����?[$�v�<���_1�9�f!/��۞����ip���Vʲc��P�X~�ƞ��>B���h�Hi�zFA� A��{g>+��?8���h/u�$,�õ�Ihg���%�)�x�1�Z��Am�Ћ���Ӹ|aT����TK�/`<��EqOjP��X���.싞��o�)�O�i�a<��hk��yO>o��К2>��')i��]��g��Ym��(�[�ygz	�����BҺ�:�|�,�擱qK�K(;i��T��P�=��b2�m!y�e���ɥt�U�WP�A��Ⱦu벬gqi���A���z�� ��P���v���{�q�����u��L�3
��wE"�����/�?h44F*>Yzf�kQ�̽�B��j�Ѽ�էA$�Q9»�q�Gɐ�I���s�5���S�|�l8� �X��旷]#u
� ��VU/�&J����0����z��<	x'�*5A��O
./Z��(�rb�	��0�{"<��`��9�وz��3"^��VH�S7&ժ�ʵ@�p�u�������>�ğq��=��%#�"����Q�ά���7�t�����UZϯFg����y~����f����f�\B2ĕ4@(�2��#�&`4W^@����?V�+�,�ʨ0�L� OEOknn�73�ɤ��2?$E<�:4�ȫ&��� �s�&:T	@cAlN�pW��>���cҿ�6|n�T��OY
��uǶQ�O��N�%�;�K1�R�Z�sE?�-����^�7�A
�
�D}�i�3=Dkp���K�������69�&��,�6�BrH�VT%'�=�e7�
=2�0	��~i|g�A�ӱ��n���S��"Q�u��{ף+�@�J��!^U����95#�,=0+��ͻ���='P}f���탟=gs����H��0�X���EE8q�����-��n��e��g�d�c&T���s$�'�z���Xի�A�o�^�/��ٗGE�f���u1
��U�Ⱥ�#���D��q�m]jV+-ۼ]b�Uc�T|���j��.���r���6��hi����O�(^�%*��X_H�(�:L耝�����E\�HZ�5�u�+�m���� 
�D�� �|�7�Q'HQ�dA�m(=s֐�d���>�9��#F�V<Lx����[z0��D����Mt?�H��g���T��&{�`5!]B�Tw`P������������I�l�%�K
���b̨� )HsX� 2��:o����7D>�"���������7v�Q�fE����z3�gO��;�FH8Y/��gz��T�ۊ�Z�.���L��B��F��d� ��.(��#�=�����H+�F��̇��_U�4��?��ˉ�ꭄJ��[�U20<���e�_F^V��������zȜ*Ek�G1��{� b2��C��NU�����Hij��W{��`��o�}�T��
x�Q�4��Hp�&�ތ��?�Iz�7:�cH9>Ӭ\Ҡ�I�
��T�:�uM����k�{��~)�t��U�4���j��1�{��8�������ؔ���Â�6�Tp?��ٚ���z<T�1u��٘$j�c%)�Z�d����I���qyK��"�ڶ�;`[�O�k�7#�qo�nJ�vh=.����%*�՜�r�x,��+��Aq�~E�a�}>�$�K3�
?B�4�u�����n�8���6η �$��x�S������Q�my�����x[:kg���꺟�U|�gH*[�,���+X���E&Y�CPCO��9�q�o+]X����Kg�><��k�'M�(0݅�
��:�WP��G/y,_d{��&��/�&�y���開��@h�yz�b��uG�t��k}d��;�n�e&��2��ǂ;��^��1�Q�d�0V���k�]�m�h�������R���	�΃o�j�3]L�8����dɸ.��v�gK�~=*?���6t��
�O�m�\�0�� 9�妺�Y��*��-O�&�\:G��Oe�u_�YZ1�hB� <����uf�������hR�kd�g�X`�T6���c����T`�YQk��9�wc�@��ֳTza��?���Ev~.s�$���ca���F���A�`��S{�:[�
x�t�pzJ�ƽ��-h%� �b�Y�JȜ��IkZ̽m��^��;D�  gH�4%��$��5Ek�b��<�a�_��������I�[.X�>��@m���ݤ�p�V�]1��/A�~�C�\�.��*��b#�Z���9E�}ihp��#Ӻĕ�rݨq]s'��prc�O���s�}67����6��ĳ]��yn�Q5A��(�`�?��,*���S���n\�9��Yt ��So=p�U�M�|?P�!Jz��n!�T�����PB�mϔ$	\���B�B�Y�5N屑d��4>��yq�S���lI���楡�伴���䬬;v]��v?0F�Wl^�1GI��0��UOh!S� l7؁���p�$)%��{)�BI�]��(#Te��I׀r�v?̘�+�O*w���-�?m8�?дL�۳A�I�u�T�U�s1��ْZ�͹)<�X�W�+�v0x�/��	g& G�\r�E��/2�
�|�.I�&��2�H�w�LI|��gG`�����ʚ)x"2 �%�F��<Kח<q1��ѡUM�&��+�˅x�i������L�-fH�n������Zi������;%Vc�㦹V�sk�,U�"M��X�>���7c薛�?��*:y%D	�U�e��F�m�v���#}}$	j���&]��4�����_U��]n��~ジ�K�rw*�{Vb��hKZ�B������&���(H�H�rHv���
ơ�0�����p`c�1���:|�i)i�l1:��uDE������x�1M*R(����l.��{����GB�o�!yݶ�I�X,~g��d*M��"@lXᮘ"�+��*7p_S�.�tp���g��J���U �����Xu�X��TLOR7�S����3�s��#�wG��w��F�j���*D�u���ot������-(�2z��+af���"�>2��K"mtגpM�����&l\4J�fܡ��X'�-|������R.�-9t7��J c
�pcj--�`D�Ԇ�t*ĉN[kWq�7�|zi�9Z'b�ݪ�����Y�R�h�J�Q���鸑������N�E<#ElE!-Q{X"�������F\%�yf����HB���qC��uÛN���4�!�+�y�E�\�I�tY(8��	 x��k��
K�S�*��IS���-�U�qq�M���/7�\�N���yŪ����ڂԠ�bT�Y{َ���8:�A8�eq��U�d�2J&(Y��$�U�/�h.�:dZ�����vW��et�Eq���^w��蕏��CJ d���$x(� ��\�����M�*�^��{�{U�+�In��חV����H��gl�� �^3ñJD"�\:��L�J�6���nB��#��إ6�Eo�ڕ���]$u�>����"�\�l�U�faצD�d9%�+fm�M�9�IF���� '̀��zr�����5�_�6x����������bU8=�H( ��}����Gc��kX���/׻����Wc���G���1�a�ԆJ��W�#��J��<��.�gP���R��gW�E�ڙ��ҁ��Wt ��DBd�G�[ͯ�� �E�ށ*S	!ᗎ"�Z��"=`�G�W���a]c� g��u���M�4+En�>ʐ�����	Rk_X�L:v�����-=� ��E�]ؘ,%������1�7Ԩ�8�!g3���7fH����s%�j	��#a��"�s�ղ�2��o�]��
K-���/~���k1�P�TBm�8�.��q�I�\�X����у�B�Y���y�)��M�j�>�J�ߖ0��q��7'2�	�Q�b������)/��|�G^"r�w��f_�n��� �>��=t��~=H�)��)$pY1cQ~"��<�ۣO���:b�`��F�'�"������ ��?�!�٢_��K�wn�Y.��
���R���9����Sg����6�����,66������G�)����^]�gU>��q!U�᝛A�d�;�p���3�-1�\���Jq��I�{1����/f��H�'�Rm���U"�9gI��8L�s`����]��X"`����n�S9���f�PT/h����rl�0G?�(2�`��\�H|F�&- д6��_ܴqOWwn�fZ�2���wČ3#�謺�WJ��yP|���	}���9���uϭ������"(�b�EG'S$��9�OgL�n�J����U�V�aK'SW=���L�h?Ax�*�U��CҫH��Y���h���e�6��{��ӟ��QN�M��)��y^3����ɂ:�'M&�!�ڵg���a��Sv���u�ԋ�� �v
���8cT�!"�Gs�.t�٩	Nz���ZG��x�+#8'ͭ�Hy�����ƞ"���`&0 ��E:ڟ	��DC0��'+�!�4��S���r����t�m{Or��[���	��$�Zנ���l][�MY:�yB��ѧ�/g}/RV���Y���6F2���޷��|c��X�gC����[Q+�ԩ�|/�X���	�:�iC)��6琬��MjPK�o�m�[8�|'"�;�*��M���c��w�������Ֆ�3�Z���y�/��W���40HQaM�y�ޱ�6��;���
��QfJ�A��U��ܓ����Y�u0�����m]%!�wC��P�u3b����ȇ>ߵ� �~�)�l�S��UE��oP��
�A�8ӷ���:�E�<hl��{i�ҳu����[� O'�TT_uy5�C��m���M_�+���~'S��͟�><H�w���n�K����Q_"c�7.�|�EY��L�D妉�����5Y���O� ����V6�Gˢc�1�	m}�#�a����q�]�|��N�s��,�����֍��q��66���)G(z7��e~��f�6�O�	=�;��l)�hf�t#h�x}��3D ���'�	��\�� �ɬ�I�{�*c�Q�"ԛ d\=e�7F"�j�#w��6���
?}dY�>�"[uM�,.�3�Mܫ�G��A䯟B	��.�>/��B���
X����D�[� 1�f{v؈#�LT:�#S�o4�P{1CV�#�	c��1ܛ�9#q�>a�E饝RǔO��]���(/V��z��(KH��zqp�a�I��ڒ;�;�f�˰�^�Y_7$��ZϽ4��!3�󫱿�P�����bIF�	"���1�g�Wn��>�8�������$�M9�'�?�݃��P�j7�3�BV��]��T�T�u���d։nF�����Ļ��h���jhv�'�x�G��Y w���df}/��%3�p��s����1� t����Yͣ�X�k�9��������cku�Pyƞp�e�Z�LX2��!�RO�����<��ٗ6f@��љj��^������K���%Ơ�c�Kz��z���#>����E���I����F��3��Z����+biv?D٧��!&3f�Ƨz"4t�<�%�<�6�K�Ո�ǉ�Ն��*sdk�W�cҙ�#�D�9R�^H���{j����{}��ӓ��rX�Pj0	��q1�}��Һ�6 =sjp�����*�l����]U����m0�utS֮4KR��r2/q���?e���*7�0Tj�A[�� }F�]e�]���[��g3�5R�,��,4WKB��8qҐ�QbN�u�*��˥��p����N� ���@��cjV�)A�J�Ot��%����� �JKa�l���؅g��K-e(���8�	�����]�Ϊ�$N�.#�V�o��b�(��X3 �A���/p��)��~I�c�-��؅4\ �(��)=&������d��]�)m���MZ��Q��P����G�U@#�h��nq�%@Ҕ��b�t���� Ne�f����h�m�N�����f�_��#yN�
���a>���:A�zw:mU�k��a���i��l˺�B��Pp��w�3�=���1a�"�ޓ�Q�ؠ��ϔ�(Dp7�z�;^�	;3H��/�����s���w�F$�P����!̫�.�}f?Q���R�����C	H�\:�s��䇇��av��e���4<���V���FBb�x_��Ӿ5���@8<'a�J�:ml�``L�c�b�h�ӵ�;S5�Z �O��01�{���@*�,]�����9��7���\�a D�M9n�jm3��7���O��d�|�sr��5�������a���sA���jF�h螴�0�\+c��Cv|��ޖ�����7�(�a_cX���ľ��+ڲ��*���p�T �E`9���-m�?`�#�Ti�(5��G����	�7@�(�0�"w���ͥx�7��×����#@ ��ntD�K�q��C�$)j"�=��Z�`�։Dm��ĭl˘����}F���)�B����4�H�
���B���IH�ae,6�����:2A��Ň�����{�0�[�YmԹ�eG�f��ϣ�	ȳ�gڊ&��P� ԋ�ן�k�2���g���K^�InH*�:�����"��|v\�s_��ߒ��%8P i>�Jf�����(��#H��A�a��t!���gQ�:ȔF�!d�w'T�b1����@��P�s2�.e�}�p3�i�ѶU�xV!����\���{\O]�0�4�x�B�bL�("@[�m�[��T7�+}V!���<�bQ��>�$9�+/B�a���]��V���Q,�W"0�;�IY;b����0=�,	�F��A��W�K��I�V�]Oi�9���q���pe33N�||��L��}ڒe��{M��t+8G�eA��.�2B���j{�f#��)���s>R^����@'�5��~�bh�Q?J�\Uc��2b�]�I�"�����	�8ơ�3����{zE�C�Ʊ6"-�ߊ�����oHk�6���X�?m�2S�x�4�/r}J0��Bh�Qj�!ݜe{�$,��p�-L�r��^�[f��R��n���t���D�o�-��j��CHG[��M�5��@bX&�i'��~��m�q�^�R1���%��)!�o��%��.lB�+��ۄ��������՜ԏ�4̬^mZ�zQ���tS��n���3�����:g�Ɇ �����ys�N��i;��2�]iz�%W�)?�&�s@v���6B�NJ�I6œ̻r�����З���ɏ�B�h�C�����6FRU�O	�ph~���{�"��n���� �R�V��w=G����,7�t����}�Oi>��4��#�
�F�E�	���SfL�1�Sr�7�+��}3+���=z�6e�z����
�G��s1׭i�A��/��۾���-�+�	�T������]��\
�jjC
w�T�o��]��,��+��)]5��{��iEc~4�d) {]���o�5+O��x��o������M՘����ǐ���'Jև&>��s��mD��O�q^��]�����rԊ�qO�&��Rc�8Nlp��QC�<g�NN�X�b�[�O�+RӶd�&\�6��Ӏqw��}׍7��}.�ŃnճkҩF�C�M�do ���4=<�<{�j?��ci(���ؗU���+Bk��T+���a=jM}�v��H���d�tuJi��X(CJ@#�p��GL,{������ɳ8u_L^{SVG]�HMl�E��4.�y�VtF������s�۸D�
�2� �8�P��[�dQ�`~PV�8�?f�&�K
ݕ٠q���-�t�]F��H`Y۞���R����S����']8���\|�q���FJ���ڮU��o��i�w�|H���Ge���)�c� ���Y&�M� ��ר9�I�h�5�������)��I9�Js�_��'�;uA�֝�ez����:�ѻɌ*��=4�:1���3_b��n��Y�����I^+��d��#��f5��e9֓T��&��6͖4id���.�		JG.���m� ��Q�"�X<���
NW{��v((���0ݏv&T�b]:q7�Cm6�2$��  ��Q\~����LFS�A��1x��o;a���9�|����W��v�-��A��@w�����x#O+�lHُ�� �XŨ��+;�$i����s�6VTO-i���:$w������{�tG�W��hl���.�eca��"�d����
C�+��"z8�h��gD>������p���)���@a�������&��- m�Y��O��H�a��b��xJ�iT�+�LZ�G&���u��ސ�(����fʢ2o���=UCNh�<^�J�����la�7�^�T�����H�ÿ�e<����*�����8�+�8Aų�LQG���D|����vy��	c�	ؘŶ�j�f+c-Ǘ���a��o1�{_�cчj��8��B�V�=|~��a6(IG���2�;��@vl����������;�P#=Q8qR����Hz0����	rl����,	l�>�@ܸ�W����n=�o�$�8`L�F���5�xp��V��wQE��w��:�ߛN�@Ħ��aY�=u�Ek���8����:$J7�&�$�mr(�.g	��a�Ƣ�˳�~��̒�B5S�rr@���Ϧ&lh "�&8�/
�F�Uv6���VV4�ϑ�Nx|hO�B�z�挑:V����i�K���]��zr�SW6}3�W���J	d^ z8����ٜ��iw�*D4�� ��P?V0e3��XV���-���k�~������/9�2۪�,�P��}��uD>��A&�zd=bV�za?���[|�6��uŮ5�07-'&@*`r��Ӱ:�dk�Hb.�IUk��I=!��iqܝ�+����n�U�L���LNxS0lo�vD���Qz���$oF�l^X�:�����ˋ)~x.�k'��f��Ңzà�\�@^���\��#����(�!(=�B��jj��Vu)���4㟂³�Һj�щB ��9&�l�!�
�	T�2 �>�Ӵy;.������Fb��9��$��T�pF�d��Z���J�#`����9hGY�����{cQ��|[�����Ƹj"4�m��� ���{)���B$mKw:QO��1ճK�G����^�g�Թ��nzf�����}�"\3�Qk2{`E�9~n]7��1ᶃ�(�5��L1���v~�׉	J�Wl��dB�&���O��~',h�r�6�3�j#���v������#L$fry;v���� 9��ڭG� 2�t��B�#́c�U�(�%w�8>�p���#>r����b�JH
��H�m��� ���k^U�����+�a%3�Z���f,�zK����ߔ_}}��/�A&X�ù�V����?"q�\�=Y<𠹍'y>����Sגu3�j�/�p�οw�Qm�2b?4�������
m��f���-U�=�0��ܸ����'���%���.
?ݫ`�w,Z�T ZQ�J�մ��t����`��I8�q��or�&�����UW	�o��_�������]��4�{{��Ppc��1]GF�6�@	�✷�f��L��P8�V��X��6��Yj�h�P	���5*�EC)7���%
lZ9�B6m��K�����M3k<��^(��\�N�%EE��OhH�c~��)yo>T���"�
>��W�~��^T�\��GOD���ݻ�)���XH��v���P�h��0w v�f�?��vb����X[���Gﴟu�oY��.dάu"��}Oj��_݊�&��D��4r�A��=���z�[[#���ށ�r: 2Z�l�:X����o�RWe�fJ�]��j{�5���W@� ���Z���mY�U�ꍫ曖�����
o4z��-jC�O
G>0,���#�/ 1>J7[f�/�61"?u���-�I�&�a��\{C�S��cS�%��^�d�A��a��A���Bnva5��2"y�&�T��y`͜�ш�C��ӳ���=�������cX\c���I�	�����֓ d89�(��d��h*鰌�\#@�r�1E�"Id�8&�{�vVd�e�����0�������^͚x0���9ֹ�&��d����������7E�h�#�Ť�2֐>��)�	@�����0��
X\��BSf��V�( �������7��r9���c�Z�J�2�z<ֵ]�s56|]�mY[��։�N��!d�Ο�%u
�V�<(�	u�>����
_;�+&���ykV�g���iz�Y����δ�:���/N�/?,�Xi���eH�a=�C���qG=v�3�h��tۄK�i�a�A'u��	`��f��ݞş,'��CjP�DP�} /�����	���N\���8�a1dN�`BΆ��o�a [�R��mZ��]e>�|�r	�a3����NƄ�I�13p��\�}?��f�8H.� ۙ:S�ub�?c�Ta�>$�5Ӎ��y���;E�㈇�8�,����i!}��Z[P�jE��,��ED>��|j f���)�9i�v�|�ǿ=���:���=�w�����S�LHiB�0yCj�]h5�e�=3���!|���$�B�^T���"������_4{�f�}{��o���H�ν�.�ShACe���w�&�Y��n��D��ڶ�xB��O([���@�����q�AD��q����@�Vۊ6,�2�vZ�U���a�����c��H��j���ެJhWXȌp5$Z�b��0�|��bJ�z�\�s�Y����t�ȯ�Ǎ}m{�4��c��?����PdR�/{��r�|tq-�d���C��J�rP
䜓�g\h;������%U�x0�;ܘ��Zگ�"�(gL�y5.���bHb3�Y�4H�%v��7�61���O�J��/����'߅N�"U��7�RЉ���E�j8�ɏB���e��~I��F8U5�ύ�9���Ybg�r5�s���Ƈ��⬫9X�p�S%�Z���#-oJ>x8��e�.�R[W��z��:b*�g쿦����3���wg �[�a�A\"��;�9����R����0$�M�V���쥵�����%a��<�+�T��{�&����e�8�&���^6-G73�[*����۪[\����v6x�#Z1�B�TC�6D3D@�׮���͜����+�dF�\���0�����"a�g	3���/i��e�i���p�!��K�5�'�s�}�,iV�G�^�g�9�*s�6�y�R.b�Ь�I̎��;�ϵ5�>������5iF����yAr ��32�2�������E�D���.��_
n�AYg��f�>�
��Ʌk_�@��� >�3�'�*�li�E^�-��e��f�4�c'��_�ϭ�mc:�S�S�������!`4�]y�{t7���~V����2fѪd��n�p�ly�N��i��]o��M��/o"�L�(���/J(I�b6!G�Oc�}��S��8�����1}�y��Z����LvL��Kr��E�_]��w ��.۱Ǌǆ����Z�ی���af�w���.-OI����S�	ɕ�0�v��/��X�t�����z�_oj��T�.�u��·i�qS�d��C��1��Q��Ì�Gť����*u���s:+'ɚH�#?{���u�l�๚��s_N(�6�ʤ��2��.���^��X���չ1�."\9����,�#a�8�+$IT���qU�^�}3J��Ί�\6���}C=�7P �@Y(��$��˰�1^�4<rKN`�[����.�>�.`\H�}��K����@�9iBx�.�=x�������y�q�[��<��<>ٴߙz�y�TԬz���� "�܇�D�hWP�7^+n�8#~��$��.���(�ڄ��t�"J����ɡ�����"��":�c��twJ�O+��}5�6H��E?��wr+�*`q-�y����_��a^p�*�),�XDs"}�3��[ij������~EU1z���WV?q������i`���'��dz��X���D���I����ޚ,�L�oz��D����OZ�q�|r��rM�!���O����4�@�1C7�I��U?KD�I�)xK���T\�ک/�G�)qݡ�pל=�Q��.�LD&��H*6�a������鉍��U�i<P��4���/�2��s%1ɴIPF��8��������eT%=n�Q�d�����+��:�CE�����c�-�v�cF���:,��7� �� ��)�~ i�l����3 6 X�+��������4���Bm"%Fo��on�r����v���"�'�_����.Ɲ�lb��_͋��\{r� ��q����6ۦ�t>��\.��7�(�<�0箊~6c��e�?���o�cS,�E�U�b�Ł��T��=��8���z�>��/-:�VTL��S���i�IBb`=�X�ߨ`4͑�c!�p�M��@u$��Tv�BQ�Y'�;�u��r1�)��|���a�s��b��ت	���rAUl��΃%@��ll*��Mp]E ��%Ć��w^a�O�F���a���ڂ.��_HP�CwS�J��s���W3 �VǙ��(���F��,�j��˞�C�G6�H�,�LpQ4��@=dכ=� ��l��@��u���&Rg�IK	-J	���ކ�k��=\���b��uu���J���A�A)������t`�Tg���
���BBs�y9y�4��T�3^�if ]��Z��$��Ϛ��O!nO��� 1so���F���PRMY�ƞ����
�h4Zn �C�S��w�������l۞�*Xb���m%`�	h#ƫS�n 3�+z8���V~,l�pF�Yc"y��6�4~r|0釙E�vs�S�iW���K�M�#�\?��jҋ��$i7��11_�%�F�pS���z��[:�|��s�h	SDv�|��q�#-K��Κ�c7��W/	����5b�y��pk��x�\P
�hެ~�2H��|���e(c�ځ2�9���^>��e54"N�~g�2�
��oC���Z��dU.��xs�5$�\�<��"�oJ5��R-��
�-�V��Y�#�P��$,翭]�K�~ﶸ�����ps������]#m��,�J�]L�Pdp5W�i�;sŝ� 
E[Lx>#�Q�Zz��IB�&��{�伿B����O"O"T���Ť2��$�HiC���z�8�H�J�Ӝ�8~������T�Ҕ�w�~��X#c�g���T�I]��`�%	9ک}Ϸ���Uh��B�c�F�w���o<3���������{���0cG���͎�=`���B�qP>����J��_r���O��TZ��v4��g�W��rn"�a�y#HI ���8��[������'�V��S:{\�](�G=�tV�g[Tn]	&�yA٩G%:T��T��[D�[���"R]��h��\�r�8*%��@�9&_���>�E��������-�N��,[�P?"�Q,P&x�S�n�n�S�M�t�$r-5��N�����U����r2����&���?�i�Y$^�(qy~�7w[�y7�!5+�tm@�3s�Ɩ���<XWɥ�=��(��ǭ:�+�}Ww�<�A������i=�l=Io�:;�w�<���� ��_{q}�%�Y��v�{$�� ܧm�MjG��	ܩc���M[Hn�&��A�ިk��v���6�b��T�W˸��]��~!z;�lc���'�1��v4����l@,v��+כ��R�(�D���c�©����e]��$'�d����/�p��P!=��i������I����-5h��b�+���UnFάsP��@0;��G����d s
��F�w����L,�@Pi�l�43|��P��㔢 �b]k>�����zY��6O�n-�"V�k�c�棑H{���d�ɴ_H�'i>�)�p�:�{�@�1���-��Y�NKL������S�����A=#iج#��)�)N��1"�&�J��<0j�Э%��jH��h-��a��ԟ�7���9�5t�X�9�5G���q[��#�hяk.�i�6����1�C��{ܑ�@�����9��i���I)���{�)�
�lo"�Y�ډ��t{��z�O&&����¦>ֲ/�ȗ�fiK��a+�`�V�v� �̡ˡ�H��O�ע���_����������v���ҹ�^����y�yTvEx̖���>(��ɷ��������0bgCdI6��{��<�U�7�L}`�Q�<�n��GYS�\D!�щ���6:�CC���&X�O�ۀ��}(�v܍M&vp��+䣾 -�A%��[)����9w�Su����Yx���݁�kx���E�����+#��~�m�w���s��x��}d�N��x��9#�����D��T2��i`q�S�=2�7֢�6�&���#]�!l��	B�n��� Oa2n.��iؗP
~�+x��ώ,e�9�ʮm�Ye6E8nSYPd@�7�7����$�a�YO������6(ʼ{��wz���W.�.�~�,M���-\ ��E0���H��ED<�|�&�;X?���R��$�:��VSd��=XK]�Y �=�5
π����8�����L5��N�����C����}�azh>ʐలW����$�ܑ�)8�I����:�,����wHǇ��R���7a��ڥF%��K��H�Ǧ
ȷ�)f�Xm�1f�i�ĉ�ث�2�"�İ7Wl��!�P�x��������ʐ�����_<�!��$ �n0n�ǖ� f�-���oRer5���8�9<���o������莖s�9�K/~�>�k�S%N��\��[����'�B�7O�$�:�z9��s[��{R�������hM2��?�9t��@S��=`� �,�����[!�e���N)t�rr����u�6������x��^��/
��jq9�Zs�{�C���tՇ;�7K�H/���0vʗҗ9�c���˦�%���}�O��ѐk.T�W�
(�
���L�wْ�"��s��|�c�Cޱ�hS ���a��MBfC�iGxj`]yRu�x� Uw��,}��I#ߎ��a�_G.<A�X�+i�cy�P�π �i�Q%C���iC�hl��c�j�JPʿˮ�����䜲]��ʧ�xe���69���4-��%j�����EM��Ec�|S��#r�� ^������i0��-n0��ءo�1Se�Gz��0�
˫%��Q��/��%��pb��L#�� \����Jw�Ud���2�YN�bZQ�H�gnc��l}����}3�[�c{r��r,ڝĶ�Hh�&���}�n,��]C��Ez���Ú��R��iX���N�}��Hңm,�=�˖����\�R����%{��ŵi��	YQ�=�R�A5������z`�IM�s.0�������*J}#�P���M� � w��)����1$M4�g�C�a�T&=p5A���c7
���3�!��4��vAxž����>�}�ms��[�6�,ތ_��x�F���-��<jN v���`s������ ]@K3�tA��B���V�g��cB�j��Si�S�es�'Pu�y����\�^2F��ENm��7����}5���z�����x-}Y��"�1(��	F��6ȁ JzH�ȯx�9^b82��a)�n*p�֐�f.��g���^�X��|(�΄]s����4a�/�],4
���Q:����*�we�Ul	8n�VG���)�%-��*�eo��پ�:������Q#�/�Wu����:�=�A�E�^(f�qB�Pev�%/�Yo���T�T����i�'�M�4�w\�]�xr�u�k ۖ~6���T���Ho��~q�>�n�d��R}�d�q]�0x���&ۘ��2�h���1�ʭz����/���8��ͧ�N�h���AEh����v�N�ωۢ,���b�1�M���V�J1tQ���}�K���Ť%����#z�
�:h��ޅ��S�׹$1A݃k�:
.�?4D����>c.�5�x9sN�f7bo?�-.*-v*̨x'*z\��W#����_5��M9�47�r��h���:_[��S�%K8/Y㎟�'����д] �Fh^�&�`)]fN�=ED����l�q���������Y����PK�S�G$����0�����8 ��n҄�×*��������7��Y�E�&�D����ɧ�_���ҲIF虖m�$�M���r�lY��1;���#�;�.ͪ7���ÆG�>%��A����rO�)_�U-��
��y\�_.�)M��|���e�,��&ܥ7��7�Q �!vy����>��ȭ����rܥ���]�ӈ�h<2?�E�r؊  ?~>��!��w~�{d�Ϡ���qBX�Ϯ:؞��`	��YBJ��/!�s�i� c�Z8�򵽊Ö��й��S���m��`I���7 �*E���j�����.�u�=�A~�Q���v���6M�T���[��d�9Q���Oe����w��[�[�-,!�x+<&�e;��X]�5��͕e &�_`1��r8�j�-c(�A�e!�	�:]ɬZ��G�a�2E���5��о|;�w�L�T	�A��4g+�:�D�@���<�9,fU�Jc#��< h�fI�8D@P@�Si&��O҉�vP�T��kG�� ��s̀T.�󬰑�D�cʕ�f%>��ڔ?�+�	C�+T�ӗR,2A��!���w�`�84�X��gy��Qf��XY���!z_�I�7 �7��@�%�@�q������|P�����]�sր͵��MOW��wO��^b�L��JdX��^�t��K�F%�%�خ��������1���R�����m�\4�Mh�g�GmIWx��U�O.T�/�g?����m�V@$9ry"�f[]�ը�������b�YB�j�����2O�A(۟܍��G���?T�{|� �y�+�P0��]�>���W��p!gQ���ur���~MJsm��Ӳ;Na���4Rc@ٮ6> �ZD���!�����xM��i{�6ɐ���Q�ޟ���1.e^w��B-J6���%�`wFZ"_4p!"���[����RE)��$d��J���ՙygC�ar�3��MNdK@��F����ցAø��mg ��Ol�]�����d��CR�^S-�k�d*Q� ׍��}�d]x�cH|.�����k�8L��[e�>�ׂ�b�-~�Q��|��,b�ҤW*�Ƹ�xY�@�,a���������0L�[�+�7k��q� �p�&�A`%r���~w޻����0���� N W҂i�=�!��%�C���Wj8� �9_<���t�ݭYz��	��B��O;�j���ۏ��{G6��:+5~��<��w�E,���AKܲ�v*P�E0����p\� ����l9�:򁸊`�tQ����I���<m�7�iL9s���5�:W�L89���b����Y�(O��_2���ͷ�$�F9�-(0�Vq�'-�G�e=�lʸ)�Lu����	1���8�o�%4��g�������zH���x��M�c�φA��,>KI{eC͡,�h�}�$v#�-�_�}�햞[D���i�6L�R\��������Ƥ�^�Ax�!(�
��mR�%�([I���zӑ����t_���e��Ĵ�G�j�ƥ �ӆ�ՠ�#K8y��`�Cm�����>iY?�=nv�=��Ly@l)����	���J�;�zE��gI��� `F�����-�?j.q�������=d�&����&��˝���Ͳ���H6R4o|{�d�fY�z���B�*�v�?M�:NX�)��`��W�{!�(^�
U;��B���$�
�~܋���.���qR��;i��T���F�~:�m�<v60�ĭ��՘e��~Ze@��Ɗ�{�!+F��~Q>�-��Q|4��BL*���s6X7�����d/@U�*I�{��������rS��vc%o���'��w�d|c��kW��&(N΃��H�煼ڻ-�XU7��pe���ꗿMNeU�9�����_��iq4bPs�&|��&)-�H��ډ)^�g��/��e,�~`)6ܐ 9�.(�d�H��I}��~Esp[��Yx6Qz�`})������̏v1�V];=��y������8��K0�̣Թ e�e� ��i
��w'~3��e�T fA֭����ۢA虷��Z0 ���)�\������y���d�Ƃ���tP{�D�0�a��ڠ-��=����t��P_����tvS�������� Ai�i;�0�u0��y�2��M<8�q�>��F(�#��I�^�Ok�M���Pr�ԃI2�c6Z�F�Md��Q�'�i�#�6���l��&]xz���y6����f�~��
�g��w���˒#a�p'A�,�4�Vs`�<)�/�ң�L��]ҹ7� ãf�՚=aH�(h���(ˋ�i2��wS����n�_Ta����S��}��uZ�\��f~.̗os�A�s/�*�P�W�G�0�� _k<���W��fq��ه��!W���|=o@G����,��������U[�<=�nwchz$�����p�׻)��Z���P6���Ѿ�6��� ��B�`.MIBm>�6�p31.�N/�a���1���q�*��xTH�L��7����v-��vd���A�Ǽ��6s���������f�{�yHܛ|3�bX�osL_3K{tB��n���Y6�-!Y�ڝ�;(����T�W;iW���XTGBVA�L��=���k�[�1W.����
���)��,�̆�܍[p�`\�t�@碁�3��F �[&d�	���텅E9�;��❵��`��K�U0�<u�}x��qh�A3�P
q�F����Y�.d�^��q���z8��w`^���c��PF,�8<�y2�/��A�b	�f�4��|Wބ@[�Ш��� �w�7*��D����D�$K_Ы�
]�����>+��EF��)r��H�1@�L���7ҿ�{?~uz8PrZ�/+�UB>:<���F"�L��BS�Ӷeg��]z#ё�L��C����8aT� �1��.�zvׄ�؆<j2�+�QJ�>I�B�뫯�������	td˥|��
]� ��&��{�9jsg��m"Q� ��N9Klk�i��li�bYc��j"���"��� �_�m]e����$5���0ɢ�J�q�e`bmPا���W)��k�r��n.�n5>W��E��R"��P�\s�YB>��Y���o�l5�(h;��ә�3�{m��iևn��$��I�`bN������?V�JT�.j����>BM'��K��y}�l�X�T�7o��E�>巢{*D�?6$�"��-������)⩝�yEP�̈�+�i�!s#��,
��a�v��֫)߁�9&�����ؐe��؆��#��Â�o����I1:'���u=�n����=��+ b��2�G<����+q� (�Ɯ��~�S������~j���%���V���r�W�%�jn�*�����Q`9���f�;�c7O�~��,}AԬ[���.��?Rr��V\:[u��}h���.݁�f rc �,4T��@u�<�G|x�fᓊ*XHȌ�6{Q�$#�Y���r��eRvsp�u���C���ŕ;�(��1;�f���3(y������C(���WO�w�N�wL��&w�EP�i�Ģ���%�Ih�4XϜ�8M����_M���mn�(�:�P�	�*=
~�Z��� gg[i�pϕ]��)�l�}p�v<'�.�k���L`w���qd^�~O|�K!+��ޙ��٫*�m�9{n�/�;�
�\9H��dCB�=�V��D_dm&���!�S��G��ҧ�!�6�t����x��,�(cO�D�w��nF�r�m�إq ["37�C����YR��O$��'ի6��WYͰd�I�p2�j^U�&�%\î0'BO��5>��������בF�G��y�rV��d����j1~~�n�B"��Te��&�R]�/1E �%��It�i���n6��c��O[����\9Q�B��Ąsܐ�;�N���a��d�$b�:_M�'���N�\Z��} ��)�c�OR^�h�H���ſ>�y\IS6 ��^R1�Xg��B����*sZ.g�do���T�A$v�	��"g����~?wy�W�<��Xs���ɻ�9ґڟ	:s�7s�}Qf�J�ú]斂kL��>�˄C@�A�J%Y�h���6H�����~�Z�H���/�������'��Ns��<�v���@�ep(�6e�C-���IU�d�H]��$����ηU���%�(:��|�A^���u�-~L3�����z٩ �ӗ|[X���;�V%�rd��}m@�e���p<��$�d0_�^ζ���]Ҫ�ӥ�q�/>�cߵ�n���-6��},��+e�����-���7�]�Ⱦk+�	��ś�_�������|7�0�>b�\X������o�oi�����u&�����>J*DR+Cq�3�gjnb�񌀁���c�}���V��޷��d[)v��uuGX��\*dLd��g���W�l4w�aw���� � ����J��j�q��Cv�5�[�-��)��O;3�{V
Q63�X!J��n��k a�����;`�>}1<M{y���'��n� V��WdQ��U,(s�L�(S�z�5����K*TE<�Z����D�*�AOC
�~��`��';�ɉ��jΧg�5�r�%�ȳ.��md�ic��6�]/{�gI��o�L`��[�*���@�cv�d�|�fE�HK��⤩�܏�p;��8�w��3�褔,5�2��!��ߍ�c=*�1sW���/]�ڏ-n�>d�y3�inDf�G|��I���>�1����rk��/�j�	cO��ʒ��-� a+	�e��A�Y6�'�eu@�Po~���?�tq���ۖ�vz�y|n4��Q�8�x�"�Lp��Po��`���&j��C66��vfb1ղ��_������9_j�Wy��eԐ�8�U(�K��z��;�J������e��>QXPL�
�X*0W؅���mԬ,�b���x�E��w