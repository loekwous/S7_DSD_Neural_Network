��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`wEO������{̛�V���؍b/&�̈́�R9ne�Z�������S��zJ����hG�f�2X��Gm�[��l\?��5%��'Q�E%�
8eRO�z
��V�NK�{⊜�b5������vc����F�(���!�U9��<�����Kg=��U��슶���RP'&�ge���nH��5����v��k����oh,���6�?
���'X^kJK>,��#���Y�l��-����2��ur�(�H��ͫ�h�d�؟��N]����Bi�Kg�PWy�79���=F�>���;��ց혷����uL��ت�N�w)u ��u��R#�_J�}�5��q�7��V�x��a(e���!����).�UI���/�������8�:�Z$+�6dV[gQx��e��E����jV��n'�����C�Iw3�R�1ˣ�tn�;�K�� �B:�����\~���.�	}����S�/�TVq�E�����0�ۆZL,�8_ ���F�
Ķѱ�6ıP[{�A3�e٨R=��k3���qfGȓ���z�0�̛���iqZ�Ԃ*��N��G��a�V��a��I�GD ����.pI�����*�^��x��
��y�=-%V,�dq�8��*��持;ԣ�>X�uq���q�,~��������AZ��]��A�3���jMtd���ڥs����1�����������S��̸\�$g����.Y�!�V-�GX�J�t\�����h���eT%��������y���$�����ח�YA^�٨
�z��1'�-<|��C ���,mԽ�*obyW�MZ�#����:����bA���i��U!��6�C��lS{qz��∃�&�=�O������@*�@1î�p�+6섇7ـ �G��,�m'��i�+e,Բ��n�*���76wB��:�$��HQBtL��$������T?N��|��j�y�����$�Q-j���4S��%��"��\i(_g�`e���
����-]ΛR�i b�С�^�(~�G-ҧ���ۈ�E��C/��|g7'��j�tzd47K�9�i��m+7D"�o����P4k�q����N3��CN),�*��]��ޥNV� ���b]��T1�#Ԑ�ju��Ѓ��ա���w���\��`yK&Dڼ�Y�޹���d���]�"f�ޝ�9#�"��d�}����	5D܁1�����Kjb�u�,0�ng:�\&fɸ�V0�AT&Z�6
���1]�h"F���@�Jp�jF�DlG��;�hw&���������b ���=J���W�6K��t�d-j*��2�r\��`"9*"a�v����7Bў� )��{�_���J.�.�s��t�se��I�^�� ��^ơ
�^;���Ӗ84f�c(�.Y?��oߺ4��Ӎ�@�jd�
?�2���q�)`���pQ늢 ��2U�;��hL[ϒ���w;ʅ��f*K��h��),��S�y"K��';��n<�+Rb�z�p�3�g�ͫ��O�a�l�;�6�xՌ�k�P�ӝé�Ѩ���w�rq-���QG������k�	�m"�p�Y.������7�Lm��1擋a,���xR�3Q"y
�`AlGs""���gL�ͼ��b��ouiC̬�9�2�Y}��3�\�c�P����M�lZ�dv��#�_E�0mv����n�|�J� �"��"L� �~���&���J��+�yZ���/
2��	�+˪ �.����Iz��-���0�T"��;��u�0g(�\���A\mT�ݵ�R
,�Ng'%nf!ga���Wx�'^��K�2�#&5m�L�K�W��҆�+�q�?𹓑e$R�G��d%�m{��DdFJ�3��YrV�9{�ר����ҵ m"j(���0�˦��W�c��B&n�:��Ǧ`�e�~Mg�uiP:e5<�6�G�-�U�K�/w�%�|^Oϰ>:�B����	߇�S.�O|V2�׭�\U����{ݓZޓ�-��,�~��4�V1�I�5�l18nF�P�����k�~�K_	�f�b'�b�b]@����W�J�}x��`�Wޮ�Ț�{g�B({�4�S��пz�#+�8B����ҍ|O���
����<BW�uf�h��"q���<J
��O*SRR��Y����Ս6�vt=oE����%.�Th��\�2J�B�UW� i����#��sŨ���A����֤��O�Mu�B;ؒ��y+C��-N��PQ	�����|P��A��G5o C�V����(�H�R*�E]w�2�/���|䅣l�nWT����/N��	}��8E4�O9���+�(� ��8$�W;��������}{�g�-l<��b�Z���#��E&���k��j⼊e��T�w�Z���oLí�C���ϋ���Lb�^O�4Y���d�w���2�{.��bt�y.���_�;��@^c���(2H:j3�522l��6�Yr�ի�T��ʖ�⽊j���d�<�R�)p�O���ZUT��ABu0�
�2��{�vaӖ���{YqsW����u3�U��9�_�o*��-�4�j��{�Ch	�MZ	%���kL-
Lq�}t� �+$h�q�1iI䷤kbY��)i�7]�D�lVE�Ǻ?�ño����n�:侵Y����5u	�%k=լ��{�Z���̬�zռA`2/���j�ӛk��IL�iFH����=K5Y�q��'.39����w�^�5[��&��$#}MB;�e)�1�=|Z#�^�=��w�ܐ5�O� ���g��#�Y��W�3�=�l�R	���%X�o���i@��j�K�.����i�P���ö�lé�J+�	���DR��;��-8�>�6U)����7/����#l��C8�ku��L�hB���Ƞ��hwQ"��9	c��,Ӳ����qq���z����TF@b�S=��|��I�.?���p+�.�Gb,bu}	Y[���9K�y��i���%zeNz��'��k�i���E]��wo�z$��U��ߊ/w�Dc�2��H��#��=�+�m�Oރ�O=+���.�.�L~��������=/7�k�g��K\d;�'ߖg��@�0��S����0H��_"��Z�G��_�>l�$ �2��||����`to��9�o�@\jN�?9�z�Q�OzWTё�u�A����)e���HB�Tz!&�2wCC�`����Y�*�枅�tO8B�2z�Ë`���i��Q�[SN���L��4��I;�nW��?�o��z-���ڧ����*0�ķ�5S���WU�ʘ��Gs�����r�R��F�*�lN3�fq>�j���'��ɇ�#����߂] ��d�q�y�펜��[���;h���[�A'�O��O8g�g�+O`���붹�g	y���\��	�X��Bi˓!���*��s-͞	�JM4�QQ]�����u)�ǚ ǍJ��3P��z�Љ�c�F�#N��K�9�?���kc��_hҸƨv���N�m��x< Z ���kc���/��HƱ�t{}r�3 �=�ڑz;��)ull�/��goU]3 �~QLP����騬q�S�q��C�K