��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`wk�~F��)t�۽�]Й��}p�á��tb��=��d�˔@[_���r4f�O��8�Ǖ�x-�TY�_��1�SWfk([�=e�UKA/���7��X�BP_� ���fT쇴f���F�IE�O�5ա���Tg��+0w*��o2���#f ��\"hk�9� �8��Ј�?��D����!�F����):(j�����Ӱ1�L�3|á<b�v�k�(e���2|g��k+b�m�JO�,����f�կp�g��ֳ��fӽIZ�A�ʰ�ϙ�J<���"��!?*g����+��J�Z��%���'���Sɓqw�}�-·2�J[xMA,�t����/H�7��$��v1�!��� �φ���^���g���(`C�0��1����d�m�>����<�r�i��#�������*�o"�#␫���I�0Ly�@R��m0�Bz�i��y?��Θ�5]�O.�V%�20`;\�/9��I���$r��%����<�YX������eaT�] �4�=<���gQ`�k�S�� Ѕ7�ʶR������m�vV�=$(p��e�uΈ�[2x�.&_�=Pw?Dy�����{]h���R	�׻f���v����sF�n7��Z`=�j���	~�>SJJKJ����`^�ݭ;�lP�	K�;���[�٤
�a�wҵO�W���n1ܗ��OΏ��3ҹ�!kZ�w�s���]�����٬!�mפ
��J��5�J�����[�����`p'���J����E�h{��u�^:�Mt��������h�Ųi:b8��1�m�]���41;8PHT�tw$W#�Z޻$c(Gsj��jG�@U�Ă�ڱ��Jfɺ8?Ɖ{���9kɋ|�ca��u���ܢT:h.�N1o� q
}�6g[Gc�G�a�j�`��HE���΄��y�6��r�eiT�Y��-��)8���1`z��(}3RcT�ӌ��
L��W$`��)�S4�:�e� un���8�]{;���΅���N���0z��AH��tC��ꁹR�ŒNeO��=n3
=k�R�@�(ab)��u6����6e�W�����g�=��`�~�N.W��Z��p�7���#�1V�"���	|���s+Lo�2fO����;c��/��R_��YA���Iʄ#{f<P���W��V@Ǌ����NJ��rto�����l�m����Ak'D�<f
*|W]o݆�#�EH�@m�wU�by�/M�FL2T�i/6����G��<����h(�R���ÌZR������r�ރ+�E�В2����nj����t������^4�n��Y�s���iG�s�x3�Ӑ�����ԶWL��c��������+vN:�b�f�C�=�v�v�9��9��:��y�-�##��;X����1��d�S��J���Lv9 ��\j�AQrz1���UTۿ	��"����<�y��w�B:�F��Cr�u����&��4ؘ���1v�k8WBS�᭓��x�� ���4�M��>�.�� ��@�Ɉ���?�+؃/*��Q�\�'@����p� �Bİ~V\���{5Z�)V�ע�����:�$~���+�o�����3��N=�TQW���ZgQ�����g�!�_�J4��_C� ��:`5�90l��q��z����f�����0PNstM����X�o5<�����������u�d�aH�w]əD�ПC�lX×�! �	���]�re��N#���aA�=wILa�VΛm�Į�������X|mA���P���[1)}B�(���Tvuԓ~���=uI=��� ?��x����PZ��
��X���ͺ�-;�)I�8�|a�ىǾ:<��s՝������b>O��6�TQ�t��]��"�?<=X:�Bf�ә�'V�4��%����K���ټx��M��[��Lv&u��c��+���0 ]�V�H ����Ԓ�׼e���E���a=v��#䄿�td�+#!�:�3�hY�Hˡ�y9��C�s�h��ٕ�U��X�ܻ���鍱�N���0������!e��ᵧ�݋T�F�^��k�����8j��X%I��A�g�ȇao���_-h��N�ܛ
C���>��`�v��,p�!4=ۢ����:9Ӑ4�z3<��n�{9�ʪ6����������+%���`�ڞ��G�u�:�|�95�7�n
�U��\S
fֿi�f����U�u%dЮ`˦��*#Xߠ�o~U�������O���'��s�fa-��l57�	s~�RL�������؄ޟ1�s|���G���W�7XwaG�|S<*����0�^���d�4��F���?a���J1�pa�,Ԉ�Z:5P�ce��$�f^�Q���`�z�5���Gس��������e�dm�yu�=R1 �3���e��<��y�΄RkadI�(���	|�����H��Ք�4�s������e�ò�Uu�?����V;,/H�T��`�W�K4��x�ԓQn�DU�Ԋ����Ik�C[���}��q�@����4-�e�O�K{Նzk��`�9ǋ�nO�qt
S���v���3i�\���ڏIΣ�\%����nP��ˌ�	�.����٧���	��[X�*go�x2��\E>�ɞ�L�؝��� ����z^��./m/�Ɖ���u���;��t�����{���3�ϺY;]0�q(ҥ�í�,�@�ߚ�׫,�`:?F�r���Mzxe/+/����2]�t�'���-\e�]I���u��q�%r�9_�7��&ڸ�O�Kb�����Z	Py�e=����ѵr�]�}��OR�������́d�E�����>�w��!�Q1 a�I]mNe���I'�\�cNSJ��-�i��(y������R���gm��N�F��Oz��eNI�Rã0o[qs�J����C'���¦��i��e���ќ�.�8��ĕk:1��?6�UuG�'w*���y*:P�']JHi��?�m��p,�_%"h���ת,�Ωh�'���w���|e�l��z�R{�\��C��'s���`��D$��;�^�}�-��9�<$��d��D���k��	�b�8k�x,=A{��$�4�5~��Y�kLdY�m�"��R�Y��$�ը�h���c�%��{�R�|�/21*u�Ʃխ�*�z�3ȳ;������+.E*��z�g�Z��s[���t���!��`�D�A�5@i��M噞�%{���P�齠u�kZ��K�4e�C]����QǗ����:_�����>�ő'tb�{6�o)h������[��IL~Sz��!���eb�
�c��BeN�1�@E���]XM��=@M�Ֆ�XS%�?d��v�9z޺3%ܫ:/N/+J�z�TK~o���l�7�g�Nl�D��~�ƀ!�06k����"B�Y�)IM��K������O42r��nlp|�u��ye��C_bn!JX �?�5�l��X��7��O���i���xUz�8J�v'v�BKrڵ
�oz�V4|��{ā:*��� 81�J[�}��jE�j������K�ި1�KH� Xg���1+ ˏ6�2��캸�ĆWL3��� �	kT�d��fv�n8�f�	��]� ���z���-`'�c�I8����	k����PA��A\���F�C {���c�UZ,>�~�4�A�#V=��ʫ�aW������;�n@��:� 
�^��B��/����jt�֓'�}��ͽ�i�Br�#�' h�!����y�G��#Aϭ��$�x��u*#����d~�Bó�]E3b� ��/�`&��=���vT��0І�f4�:a<�!�wD����a0�m��a�[4f�˸�>Lh"
z8�siZ��ϔQ6v�p���܄���H:=1C��R��SJ�2g	wH�!`�D�\k&�ݏi����$a	�F����{��/�݇��S�|���,
��݅b���k�WIy��\@����$�PAw����V+�V�����{[xweb�V���1�+�|,��9�QȊ̇�疔�Hh�'̀�s��;�b��ag�����w��F7C$�����mCx"�D*�&uH�T�W&a�L��JceipUu�a�)�!����[z�z��;dN�C��H9�"H�atS�%m� | a�~��e�!�x���� cI{t���D��@��ϧSf�l�g}<e(��ӿ���+D��_{&�������($�/hS�ny��FY��D�D1[ԕu���������Y�5��`�����L�g@#�_��o.�G�o,.rN����.��q}�7^WHRf���4s��F�O)Zhp��ΧX�T��1n߿�aC�ܳ]��u)��}84�C<e���;��mE���׫U\��B�.�#0���Z^@\���H�^���`��E���c���	��8�$�4��]��,�?Ό��6��ԲN�v���u����ZT4�^t�e����Ʀ{�����w���M�~�ai\t?�K���[�W�r��̴H>�ŰYXb�:��l!�����_~��hU~�/,h��9��R-Ӂ*�S��e�Vu� �`�C��ijm�<\��{�?��V0�"WR��߱<�����x���4����$AQD;��Hv����i�p�X��T���o:�@|B���UD�5�� MC ��x+�,�w@x~ϋ���:�P����z`�p�|75G��1;,���IR��j��j>��ccՔ�[8Ӣ�L�Pr�kN�\B�HO�Pf�ƃq���ጪlny��GY;�Ў���$� 	
��|��%BF��	M����U�*�}p���̶>7��f��^BP�{��x�a[*�o��<D�玍�l��
�0P������#��׭m�H��N���F\�W�w�;�\��b�8�|m�0q|�F����L�v��9#���	UL"�6�J��c��@P��q�ek7���"�byUtN�'x�GEW����z!� �L�?L�gTP�h��ñǾk04R#[�A�>9W�|������ҏT��2��$(*\$�:f���B��ᇣ��TT�L��Q�3��1��4��}��91�p�Ŷv|�j� 0�}�V,!�G��H^��7y#*Hy��B4V��F��+����u )�𑾆����D/��\O����e��U���2�H�Mƫ�B��z4S��YbS1J�U0�#��^PQ̫Yy�%%B �f���-~~Is3��f͍8�V���f�bjy��M���9�Q����.Л6�z.�ƀ��D���>:&��i��������/�k��~jW�:���9?n��D���י�B��w=u�L���F,w ,ӈ�񄀇"eP���1����I�~,I��PVW���B���k�F����+�L��-����Q� ��W�86��&����R��!��]e��� 71z��N��Į�V���su4�Tg���;v�,89�4M.>a]�Kz&ʝ��b��`l�G��N��
j׿��e��m��IA��;v���z4�z+�M����q,ld�tL޽3%��,�2)Y�0>eu�#`�`߁
�,�����)K��|�����1t��X�?e%տ�BM꘡�"^���4LBy��=X6K��<O0LR�	E��x��)��3#�O�<LMO�"�8��Y�rx�@�3I�A�Oe���]�̙�1�#ˑ���,��nJ�d��D������f��ֆ>P9+$U�˃2ZƘ��L]G:M���i�t���D:�	������Z7�` �g�/��
P-&�{e��'��
��J�jD�sFD3��M����l����/��s6۳"��^;,���eu��$�b�L����pc�b�흴R-7f����c��� d�}�)`��+��Qo�Cc���ȃ�cu�X��w}^�BS���=�eK����>�w��2^5��Yp�?�6�9�4�z���>����������L�����<^r��L�Ҕ$� �?2��rN��A^���2����,�o�3���e��	��T[�K.Z�^��F.k���1hibozA�>)xW%#��0ו~��x9s�ھgSbm����Ta�K�.�&�J��A����żɟ�ո��R&��t.�	d+~�s�as��q��s��:���)���Ԥ��y�{�!'��nGo��𠈐t���b�V���z��-n���q��o��B�#PX��b;����Ҫb��Z4[�\�{�+���T?���)����<�^��v��Ӎ��s�I敭q�H�V�#�L��=am{�lT嵀�UH�TE_����;TKZyOI��8E�·I�҆<>�MI�B���ګ��l�w�Ejf�wQQ�{s[L���`O�ƿP�m�E��yѧpG�A\��,�%���c#/�n�
e�>[�|�bS�wG�a7��U-v:˂mR��U���J�`��F��������4��_P_�2u��Cg���M?K�����n���n}��)�=����ٮ[��8�)�����a�G���a�k��^�% ����4�FF�l ����M��9b���FT/Z�������iB�F���r�K�}�y��JrP�/k���b���H��7��m�pU�'�0o�����HL�x\�<��� �V�E�6���xs��+t/��8���a_�2�/�f�s{N����F@�q?�YJNf���R|jVb�D�{�5�|Y�_���zbn��c0��Gp^ϰ� ���� "��pX4rrN4l���e,���ك��;Zw:�.z��^*D+#N��������g�����-���h��}�R��J.�� ���ߨ�c�S�o��J�(a,��8$e;{�<�_}�i���Y�C`q�lx�3\O����3��S%?� ���o_�]�*no69<��#�[�%D��0�&ee�nQ���B�C���|����KIG�J��Y��hd�p@��w�������F���O/�on�"������V���?�P;�}�VtU[&���GO�+��R��B�|����Jb-ZC�]�ʻ�J�>����޿���5����l�D�ԥ1�BDW�T'_��_i�j%x�+��?q�FQ�	3&�,&��Yl�zSn�}1�J�~GS�F�F��D�5��U�]��,�Jn�J2%�չם!TܾX���=Ъ}޲�dXWh[E8<��'�������I�(�����FT�M�P��>��k��\@/Ԓ;g|u��������^�q��Qe�Q��e/7���*����e7�o��B]Ge�.���r����B��������%�C"��%]p�qa�TY��!51藸yo�f����S��������'X�<^�u�vȱ�'�MtmES:q��q �+�@��G�G���A��#��Y.%]�v��u)�a��l"�Qԁ$�3�����7%s�w� �S�vR��]\(XB��c�;��<�c��tpd��ߞ�����ch��3�BK3��Y2)��s*���İmV)���=��8p�W�ܙ�Bg�ɿvڊ\F�*6�~���8\|���#`&ͬ�l�^�c���'�Nf���$���~���m���;�nk���ȖY
��EZ~���\�G��RH�֟�@�I�i���c")��v��*����j��N��t���x{��* $�hqG$U7`9}�3I�o6\�����tc?������3�R6ٷB�������B��-)��<���`��Q�J�n��њ�����<���G蜇 ���y�������MYҔ C��v �j��Y�$'�#d�B3Y����.e�8b���'���?�?�qQ\�2`�ϔy��z��c�#���Q�u�v�F%�z�������v_V�I��c�pt:�bA����xy5 ~To�[��~��9�ω�a���Ӄ]~4�Wn��N�&TCJ��rޅ����M�l��x�n�Y��0ǘ��'��T��WӃ��6OY�c�̳��exjq�rZ���Қ��Nz�P��X%�����u��A����KX�Zx����;�e�(s|=��&�*�T��̑7����ߋ���eZJv�G���"2
������|���o�z���+�,Y�F��[��q�c+��:��]���S���92�|g�����$�&��7�(}�ԁy�^0I	`�P�W��Y���bT|�T�8���^5���Q�����G�#k��1>�*ME�X���s�_�K���dR��������h;��ַ�'��;2�/�,����E	��{�~1�&�Uq�y����ܚi��LP�D���D�����~���A���L9ӏɈ+0?2��$�
Pi`��u��[Aخ|����\f�1W�P��G���t�~WC0i柃�{�a��0�~*����W��1w�޸I<Cz���F�9�	��)G1y��`}����9h�iM	����Fƍ\*M�1"w��p�>k��);��������'�GQ�����&�����:DMi�T���&��%׹�_�EYٗ>Ug+e>�	~��	��̔Z�g"%l�7]��0M�4��Ix<�����p��=�z���d��q�8q�{�����3"@�u$��mk�U���`9$K���bd���Nu���e��↌ɠ����o��6�S�qk�ˑ*Ker�����s|6j���R��W�1�pmo+�5�7�+�Z��c�S��˩.a*�(H�>H�J%P��2¨��P<E�qǋ}��?�Ѭg��zHaP.�� ����/<ć�R��n��k,D[3N�'5d���"_V)�/�?ׁ=��o�_�M(�=t.��Qn�V�����L��/��3�=N�w��^ACS��/�]�},u��ń��-�����x�N�pˆ�XTN!\W:�{�G�OjƤV� ���'S�h��k�\n���氍R�g��~���)���K�Ǻ�=��L������$��h������ʨ�Z����\��iIn�-�m8.K.��^U��"j�N�7����n�^A��X�θHU{)���,;�RۜH�Q�9�7�xڑ�l�=�"�ڌ<b(fQ*�����#�k4^9�[)ϷVfʠn���Ѽ~<�S���NR��).��� �F�m�b����%�1��N�Ev�>Ȗ)�3`�ff���,ʼ���P�����0�M��˛�L��^�q�BF�� 䯼b�x����Ar}_��Ǚ���'�"��O�JWN}K#�)o�WR� ��[w��#2�̝h۽��P'F��s�*�ݶ�>�O�$���ֶ��Vx4�c0=�,Pgl6���I�1��$BԴ���u�@�Z[_�x;R`xWUG��A�`�z��0D�O����{9�E�SdV��4_�x�H��9��܂Q;�7��0�� �>FG�譆~Qt�
l�zy��hD��G]�4b�7�]F�j�\��$ez����n.{�p�o�j@KJ�:���i[P���ɩ+����ikl��(@={���}����4v/����>�E�ݏ[_=�?���g��7�(� �e&��1*���Fn^&���]��(an����+Q9�ǚ���`�c�k���P�;����`�j�C�*��O�v�t���;4 j������N?m����P�>�����c����xحxe��MڴSB���Z���	�TE���;�ͩ�ѳpn�]�v_ocN0� b�X�nFGo���v�n:�`�Ψeaȡ�Xi�  C�t-��-7��L �x3Z�5��@x�;��ZZ������pn�+X�f3�V�~����Q�|a1'.y�>����8П�!a���b��wTRX�+|�ux{��!�J�{�'&��S���� j�H��ַ�o�>�r�j��vs����u�3�2��4&K}Ӆ��j�N1u��c��b���(���v�r�_� S\c��x�S���S�����2�	T]W����4�&,&D�v9�8�
ђd��#b�$�?ð�Pb�w���/�j
���Ļ�	�_?�Ł��
*��X��q{����2&:ߔݰO���w��*&�WIM��YMp$�]�	�_L6�OȊ��R��:�Ĵ9�-��)Ϝ;^���;��b���K�zH.�S�Z��x����g�*���L4xf�?�fOu+�}S�5
n^��B�_��k2e˷�.�J��+��&�9<B0CA˶�����Z��'��E�!�Ni�ʷp_�6��
��$ɂ�⁇���*5�d�����(?D.^B�*�Ϯ`��D���}��ZR*�ʦ��=�+��G������MH�@K����$m<�*"��:��1Q���z3�R�� �^�I��?���5kHau��DQy�^��H���<U�|�n{P%�YU�?e�EQV?�}%fɥ��B&>?ީ"�AC[߉�Ɠj���ÏݰPF�����5%��,xX|)+��ԓ�=��4m�T�ζ��\�
yղB���U'�^��2�9������o;�v/����\V�#Z����BY����-iċv.�2��8ՊVB�׊ט��Ǒ=�i��}���'����<�'㷰I�K���G�l�&�$���<g@�HC(���]��~�OW�4�؎����FN����)���n>6a_;e�X`���/����|Æ#���>�&N�^^Bn�m�����ö+��O�,����[:�Xr}	X�\���ɾ�U�:8Z�l�
�l!gՋe���`��]���bjm}9�=3�R��	�F$8�y:�Z�W������2O{�!����� x^��11Ӭ��N�J5��o��Fa�t��34;���~��o��u5����/κ�%��j�Ŷ�^��ip71t�RD5�I!�W�A26�1^��.Ah�Q�~��>� ���1�SKu|1>����4��F���Fp��5f��)�����ޞ�;��]-ȫ��Ќ�WJgm	��g��{ݗ����[ U���M��*S�)���[�ħiTԾ�h,�!� ��	���.ښ+�i���}HUv�K��~|���Nҭ��$���A��FLA�uW�Y6��+]pU!���>�d���8��=�F��%�)��M �3���O���v�ҍY�L8���)K������lh$������8�#��-�D(��4��EHcH���]s�Hl��"Z�̱�i�ԯ�tw�3�XWQO!dĀ��[��}�H�"M��p�
PT���	
�ihC2Vpd5j8ث$ط�Ƌ[�}��m�Y��
�sf�qߘ�&|^K�~��O�R�-�b����8[R�p>w�z� 󮩐� ���'_�x��|c����U�됖td�{ؿE�� ���=#�M�3���L��� ��6�g8�fs ���G*��V��۟8���H;�q����B��$Z ��cGxn�H\ ��[��Ų �˲W���	�"��Z����!Ws�3`���/�b�OWd��l$^A�����pt�o��c\_i��]%�p9þ���F A�o]
e����R��a���7�+Ӽ���5�0P�I��n�e/����m�\��:�| ;h�|}f��!�sIL��P���ի�\��>�� ���^j"B��l���˒+ʾ�h�^&C_�c�4�p��Lq��+:x���3\Z��
�g���X��*V_/�.n,�4N��|<�?��uN��M�uy4��X��6sJ.��t��ܱ*�r�9>�`�?:�L䔁H2?9�T�a�E���R^Wt�N���8�.u�ֿRRd,���nAD+E�	}I��#Y�>9��W���&j%�!:V,PU_d�>?h�L��\��������VE2s��NF����|��Ό��H��l��B�􇿾'���1I5���S,��Ϲ#^tg�~E��/͟�Kg��5.��4��c�� l�d�@��>L�u<�J:r��ߛB�.-6�53�l���i����8b3���(����g���R���_�b3fp�H�3�F��.��v��l���m��v5s�P�}��t����l6k���%����vv�z
]�}8'�����Q\3��\'�|�_��ˀ��^�i#�s{[+�V�+A�VmE�NN���7Q�b��bGʭ�� X�҃ {_ju��B$W!N�/���?��Z���X9}�	�?�v�U��� �2+��]1Q2x�ɛ����;t���&:�������z4�~���3/9��j%��?G�ɇ�b]B�Q �.�P���邥*cw�N1�S;��F�nq����x�� LĜ��7��E�6���;�����Y�2A����_�*	2`�{ǨH9k$��/��FtF�;H?���>O��U���MB]ђ�?V�f�2Q���"o# F"��25�j������f3��1~��T����dXT���)��M �J�_�CLi=�2h���@`q>�`�S 9�<�_��q_��/�����MY�?���x�����2�"Ki�&��1�$㬉w�����X��+`�g����4ux�dɛC6��
����l�3'�1p"\��f亁�/B$�_�2�������*��E��9q���u����j� lxRd+?�� qNm^tp`l��PG�0��d���ƶec��*�,�������Riݣ���� r�<��{�ZI�pп�%S�m��i5�jK+�cl���	�)���ܒ�SDKb]6��~�mW>�9�{�KC��:�[�sh9�q`Ӎ�d���|м�0�f��@N{j��JY=��D�Q�J��,�� p=*�iA]sD���w"�[.�5�U��"|��MC���J��� ?�+�R}�p�+��A0�V!��}+��n@j���;�K����*��|�����>����k�Йg���c+�W�e� ���|j�ߔ���d]�XH�k�a@p��F��pD 0��I��8l��_�cv�nj��������ϟ�|��FP��Q�/��dO�����!U��(�9a`��Ҍ����6���t>�Cڎ��XS���rkY���8��t<�gʢ4p],����ื����>�Eˤ^���������b���"s�1�����
yu.e���	��o��+���%\������/�囷�d��{����oC�a@4���"w���W�U�_��f�E:��d"�0���Re'��xrtgA�p:���Q@O�ڡ���PX�#�ԁt��&��q���������J<�N��x~�V���LN�\��kV���WmGP���eҰ��������V�N�d�"{�k�
ʊ2-�~{K�ۃ�N%'>̧�틱#ޑ�3J-pw�p���\�w�
*N@�@e��*a����l¡R�;�&���@���l3f�
����Σ)�~�x2^|�\��k�+���>9H��! [ds O׮�v9���V��/E��h��/'�D��ɮ��]��e�B[���K�����U7��}Hϐ���������V����fRٴ�RS;�q��9p�&�X�l�ư��	���K�k�r�19&���Эn��fTܺ)�_8�������������:G�,1$(>پ��?���XJ϶k�+�'�(d�V���5��|�^�i���Z�rJJ��C�p"�a�l���i�:o�j�K9�`�����F�;�"��`e��B��Cm*��"�+
xk�4#�s�a�E�Br�p���w�՛������O�Ji&X�<����P��Wa`2��)���9��Խy���Y=���	���;��l#&q�iIa\!��$��쑉sx`�����!@�6	!7�F�V��gZ���奫�5E������gD�Q_u.��*�X��/#��Y�9�5����R|7=4�7��	�6�q��;D�EF��*�+��gf���� �f�� /t�S��hu�56�%�(A�)��N�H0�����h�W6$
��78j��E���/v�e���9M^U��*t���K���7�'��x��=CQ�����8�e3s��j��޹��}̘���gg�~q�t�p*M��wƘDCco�X��c-�Y\>�u������~d�"�nc7b��5�,>�4�[��T��E`�$%<���G <��a����V��ct�{8�lK�aP[ �����pl�-��q��,�ܷ�jǺ���rҗ�B�:(�x&��i�@υc���_�Vc�86P5�����@�%`hew�����m~V�(�x�[$#���'`��\�v[&lI���\���#��)Hj���M��)v�H!�)��C���t�_�FM�!���*Q���"�6�E�䏌�bb�$���Գ�_�Քf"�z��(kh��; Z�i|�B���RI��0��q!��֕�=�аR�����ξ�@7�P�D(+z��C���OE'DI�dL��"�kS>�N!�md���Ze�?�W�s���_)���� >j7%�0���e:���Ib�M��ud���mC������d�|D&���i�:E�R��?�ټ�^� �.ƒ?����`}c�����}՞�hP�u��A����4�� x�JFR"�A�X������@Z�s��|�R����M��ȳe�[��1�M���/kpPd]���*�4nMj��ų$w$2^n�*;p����2ؤ��t\�u���4��U��DT���%׊�K�1��<�8�YR���@+m�Ƹ�h��G�1	"J��V/��%�S�fnQ�/�#͡.@������s�/����� �ј�7���r�`p;
-��ҵ|ݗd��Z�C��@{
îr�*�z��w~�P�=�܌D��<��<���{_g�I0�*��POn_+�Ŧ�S%q��>9v%i�<�vYx��X�n�@Dê�]�B�9x~{��HBQ{/�T�@5�K8)�Rs(���<%F�ֿ��V��8�W��F�n�����A+t�쨄�7fĵcj��z�n�D	��r�2�F�t�W��/�O%2C�7�b͐��wP�y�hKV�2�o��Y�&XP:	ل�ev�Cm���s��i�m�x\|C��(7�Hc�z-7\��J=�V��Ϋh�T�z��Da��BUNٍ��w珉�?��ͥ�_XK��X��DX�@�dW���//�݋c�X�v? \y�f%[24����_$������^l�w�����D���%'n)-d�g�%"��Q���2sӵ��6�����6�Sߩ�w�y��TQ@k��;�m�����=�{��=��^���g�7�V}�����	m�t���Z�4q��0��A�k0���ٶ�R�l��X��y�pz��!��*6Iu��)K#8w���)��I��Kym`n��d�;�U�����S������աʊ�_Ny��R��
��b�]a'���pyP:].�1�nه�}m�/1S�QE砋�t)�E�s���[4Ӑ��F6!7B)�A֌;�z2_�.���rg�8��[kˊ�O�X`�,�p����$*_��V.nK[P���ҋ����S��l��=����6q���ШV@a1�X��L7B1/��U	Y�q�8�����RQD�ǁs�Գ�+.;9�VH��k<&��z�HW=����
�_%ǎ���}��D�!J����uY��/Y�5��V��D����p�'���c"?���p��"N������L�T�"ٳ����*���b��FT*D/�b�(y}ٺ\�Xy�_� �T�e�{������@�V���]�_)�l�CK�C�\֒���g�3���vSH"�ܰ��K�!����R�}�O���M�;�|'Ն��>����NO��
��0���ez�2�����3VZ^Y���D4��pI�=�	9�0�~�b �-go�DX��z:8-U��B���`1�PT�9��9����GKY�v��_��5m���ϬOc��mX�g@m�������nQg��^�Gٙn�ޚUXU�4*���(�ӿ_�!�N���]���^����A{�R<1�	�sG�G�Nw�sY�)a�7}���?��m�GYO9~����y�}2�%Ԥ��$gv�d+�kc���fB� ��2��i!�$�p��G�:�ը&ce)PF|�nԻ�|�Q��`��I���!yZ�l#*yi'c��7�~�$�z(��<�(�x^���x��m���$|��^@����^G����
g�^f��ȋ��&|M��1��B7�:oȿ:<�L�ú��)�}��̭���Vb��I��w'� �A�8ҩ���KY����T�)_;^i}�Pm!��ݘ�r>*���;}�%�c!�+1�
'9�MT�B �{V5���_�ȱ����h�?(��}&�#Uq��|}o�i��7�_Ml�j�#�s7�"��^+�[�|�Wm8�6~:������&.�׏� �ݫi��:Ox�q�W���T��6��;&f�D
�啎\��8�vl*���4���{�+7�����HO.�(�G�U����@�0`��l�3�Ԑ"�hd�O7���!�Q�*m�Q$y.���5w���vP��Jݛ����
;F]�  .;=��:Y�T6��Uvi<C\7v����R��MH4ĽH��v�W��`����TwB�����ΒQ�6�/�Q�4	�U°CL����A�P�v��B���� 9FBN��Ξ���8�'Rc*��t�2-��=��iGcPY0�>}%�N��D[@�j@�ې�� ��C�vu�f�~-�AN	��������Bض�q��>4�cs��"�?�r�=�F�����,?��UR���~���|����1WID�d�Zר�n�Sj~�uB�sf�^X�u�	 Y�W$�S�+��U�W�<=3�.C���� <H���I�;�`�Hs8�i���s��q >�w��"+��*��V�m}�u0U�GIU�<�00�ѓ~�\��{�?�TmӾ;(�A�L�E�+#��֏�� �)��DG�U[�<�^��.b�i���)}���|�&��;�yf���JV&-Ҳ�j`?�7u�=�F��s����%��(9������,�ݴ{ cUv���|�}q*;�7D[2���	��l�V	*6v��{���� �
�FN7���ў�oڕˬיWs�ەo�J�`�h��IqRM���Z7����w�i�Qƒ�4�U��C�+�[{=E�2�5T�w�I��#���~�<��>�`���g�e��r^��ު9�E���T=��4L�INµ�
7$�͠f�nӰA�ɓ�Op��,��5`��T�k��mc��&C����բ��k������A���C��� �\C����.@Р�5$�� �����Æ�0�v���{�,*g��,X�����ԸJ��Z��߰{��_J�֒�TI�w����}F�<Z�d�v�Z٪�5��=�'h�Bl
鋉��nB�T(a����ǒ�*U�MiLN]��`�������Ō8�V�~k]�oyc0@As�G�O+Wm�%����d!E���5��a��1����y�w�P�C��r��&�GK{Z�� �[�5s0��w�II`�w�'j��F[�ļqH/�mv���5��d�$���t7�ϗ
Ph}�xd�RD6%���̾5}�����m/P�,MA��[V�֞L���h��l��J�HK��ᔎ��5ݘ�G�o�C������7+��HL�8q0x��O�ڦ�+�qXCY��W6NA ���{�)�F��H�{�n�.S�%\�c�
�W�j����u��]�41~\��qRi����2(�y�Z�ZB{�A;b?@��,a���Z/ABg�JjMr)����/��D�����wR�}Z�}lߖ��d$%�?�O(Xa�,���ڶ��m�m3[.����"����~;���N�������0�L�`\�I���O崔�1џ��@��jK�K�0�k;O��J�����ݖw4�B�/� �P4�F�$�+Jj^�K*D3�C��_�\��-��{�KM������n�Lʠ��v�-��e��&\��V�+�T������m�s }"gY�Tc���I�r���P"z��Y��_�\P .�~�]ws/r��V],P&�  �h:ߜ�;��Ӱ$�&�8���.6�~v]�z�a��D�}(M�G�fƩt��L�WW�/���8�i������,��c��'�_ҤV�٩{ ���#��A��j��j�$��X�j�~cS݀S#�i&�i1����E�-_��ؠ��hL���/�ȡ�o���D���Po|������n�w��vF��q<��C����D��4>^�Y��@�`n��Av&MЮ�'	���i��s���jt�#����Gp=�]��7Wj����pTnE�b�nA�Y=^���&Q��^��R����> �C�.A�a���}	��/�_�]zC!�H�QBՑp����tt#��o�LV�h$�:d��	�07ͨs�<p�X���=x��nՓ	�L#�9�C��Q����m���� -��-??��W�@x��8pTY�d\f�1�y����� J�/�Ú�9�M���У/���Y���K������S�|�xbE� ��.�^c:X-�H�\�Q�����
7���d�ϑanϷ�$����5�!�OAߨ���T#�����C�`����x�Y��U�׫�^ �Ę����,�S�v�]f���JĘ�@HX�8E��[��z��+��� �X��(��	�L�f�(�|18�A�_����Q8�@��5��-�gVU5����E��2����5�Gq[�!¡:�\�����m]6����:�y�v�!��W.߆�Xm����a�,R�d�o�P��ҁ+�d��(�����`��+Ԩ�ߺ\ڎ�8 ����=�-��b���gOc���q����zi��;V����%����ԭ�lc���Fy�o�'̞��e� P�:c��T�T��"b�D�߻"�O��/U��"�ee���隋U��	��q\��qٞm�v�M���[���ry��וg���"gt�=6r���׽�EBQ�G ��g[qV���ܯ��7o
m����S#ƈ2s6���fpa8l��ңr1�i��?C���Vk��"������K���z��HB���̧H���AŁ(�ހ�A�;y�m�# ����(+x&�:��@��o)����ԶW:U��s��m�������9�-8�EQ����Wt��)e}�p;�)`=��_��U�O�7.��/�o�V� ���=kҚ����`	Z����V�PR@�T�Z�nw42m��O犉ܞ1�yK�39 ���� >�jӟ
���VF(d[�E�$B?М��, (b�:�3ӄB0y� ��tJΟ���%>�s�|��[�ˡܑ�`�\�4k�.p�[�W������9��%#+�	�����g3��������{b���*���c�b	ܷ�P�̆�S�Б��Z:��2"�����ic���]�����������^�	���=�1�n���t���#Yy/���'�gD�]}9* ��J����e�Dr�z3
���C�WF�{ze���xf"�~3�~i��lX��*̃<<ӑ��{`��3)��ϯv\�r��x����s�-����#��ړ��V���.��'Y��Ffz���b�KaK\/�`�B���I�-�2?�F����®:,
���'h���,9Z}�>C�x>A[���y�rV?p��x�.B'���.s��cG���Z��Ex��8ɪ�(��x�F*��q��:��u����'�K�"%V4i�uL����Wor� ��p�$� [���#r�����8t��uGa�N�k͘�ǦϿ���vU0mG&�3տ`�k! ��@%Ec�C/~�|����&z�s��]����N�L%�v�M��kj|��o/]�|#`��HZ�nW�ؒA����	�!�2�ABHI����J!���e;�\����s�i�1���H��@#K���g�xk���b�q��-�	�1��*�QT���cy�p��DF,��������D~��s}��n�Ni:*{�2��t�+k�5�j6��`��^ƚL���0bWM� t�A�HB��C��lk�;�Jߐ :�&��#uB{�"�z�������!a���/��_�p��CI�H��i���n'�>&�ـ���D�ڏ���XV�3V�n0�C�xfb�\���bp��4R$����ub?��~~�6�G\I���z+G8w��Fm�� 9�Z��W�����Fó�n��:-���Cn��8��,sxƛu2��d1��!9�x֑ ���������j�J�<e�tc�{$�{߀�6��$������Ñ��=�?η�|�碋��=]���(�7��s�U���_L�7���!T ������cq�:{�~H� ���{�s��"���n��]'X�Ń�d40�<F��G���y�EZ��z���&��ן�z��a�i���N7/^rA�U]���4�z���=��M�:xG�2�>�_�l_P�3P���p'=���A�~0�.o�x�Mu8˂��2r��zoȺ�%d��B(=�LzP�(k��:��ux)���׼����"����Eswӓڜ917XՏ���.���ˎp��Se�n���"4�����P5���QDI1���WT�o�EԾO	j����~ܜ*�A�vW7��%~.������f��.��V����U�r��s�K�.��><��Ǡ�(H�;#����ş� ���<qo���Vk�"����T�Y-c�;)_�4��2=�)���rQ���Vw5CXt��s,*��K�v��s��.t�ϧpB�V��(���V?b�f�:�G<�O�P��xB����ܥ\b��~.h2�e� S!X3\ئ=v�}�E(�����J��#����IF����/�~d�9Fh�D;5�w�]^�5<=���փ���9�Kҩ�],��p�.tӛj&�L pu�yǵ���cਖ��s�:?G���U��K����l�E}�i�-Hh��g�Gd�5���=�Z��l4	����x��̅�*��U��-�-��E�5�z�5��]Ɵ
0��������}�����~���D���������Ú�J�
��f�>u�.��K�=�)&�u��s �ؚ΢�t���j�N:sn��+�J��㲄��K�f�Q��֯{�]���8����/<�Kz���^���F$�ؘ���W�����qI�]�9����g�ی�ki�{$<���9L�Q~�=���w�ı~M]�
�o��`Jf��Q~T:��*?��{0�7݅����6ՁX� R�Z��m �WQ�R��qf�m�01�y��U