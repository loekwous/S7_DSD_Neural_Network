��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W����(t�c�
�0���ڷ��*D�]ׄ�vz�Z�k�,�G�������R/i��S9���Ȱ�_;B�H����R�RPP��b��� ۩���?�lв��t�j��ֶ�=�?F�A���{��?`-߸���I�I:�L����\��{���R6����k��j�"��lg��-�A�,h8�O��9K� `�RDS� Y��Sl��_��0�ˋI�8*�m-�쫮0e���MBSz�O�nW�#m����zq�O!�9祴f�_Va�Ht�}�O����g�?�p��p��V�qi��R
j�A�j�_R��F�b�O�Q���?&uHN���^���撉ց��]�뮪��o��;4��߄+�[��C�>q�c`��H|jX����]*�EA�1&���ғ�WD��L
��̦�����h�']��f7M4��J$0� _��8w��!�y����M����a�3��RZQ�y�S~N��N�yzBSA�_"�?)Q(���yf��P"Գ��1vGB�%!hlʝY%�H) b��4�`�z�i,�K��5oHR�|�����0���Y�E�N����;��h�v/�g&���z=�R>��I��m�ъ��MZr�/k�e�4.�f61BF�@W�F�Wxc��^�x�|�?�&ɑw�CKy
A 
���'}��`18�S}u�&il�g a����Pv�m�-iS�`]Q������{�9����7�d�5�׶ܭ+���[���>��\��������t1���O�F��'V���3g�h$��c_e�~%��iα 1Q�	>D��?��=})��\�����M��/�Wﵥ��<q�Z�:�#�!=-9�lޘ�i7A8����I��r`8X�vN���[I���03~��[�Z�|L9&��J��G�+>���C�*M�H��q��i�pJ�-w��HBp��P�J����3����C h9Њ5���V�7_()�~T�TBH~g�ˬYqeנ5�����-V�Z��Y���J��]�K�.�^�k�O�m�q���������ǔ�f�Z9�W��ޣ%�0�ܳ�W��JR;E��e���ߕ����
�f!^����y+
;9�1~��'-n�kg�T+ג�� ��-�%�L�*�p�TոS� v��#�4_����X.��J�@]��$&�������I��DN����wyn�A0`�zu� 3�p�T���qJqq��� א���=�k�� ���|��0V�s�Z�� �5��|��&��i)��L�h
]F�u��$�����A��;6�Hh�ʅ-�m� ��e�)�� �&��^O�4.	'W�U���O%�X*�PH�*(���ƞgi���u��p̾�N|��e��0uha���&5�6�*N�cX����N� yK�J��2��M-�j�C7$םA�wOK�W�$��vdJ�M��զ�!H�� ��	G�K�����b=�X�d�`b�ʾC����H �Kv>��[�Ҁ�*����m�ء�������� �l��x;�Cd�U��yǄ�=Ic0�\A�-c:��|���L��̴w,����M��ǿ��y�ǟ�O��Co�/�g텿A�>a�O+���k�;u�6w?�o#�|t�����(�t��:zH�G�A}#C�����+rfB��x���U�½/�m�S��~<O��;��b��i��g]W��yvE�0�+�S�ə���p���H� J����OӦ���0���s��o�L����r6�)���
��G�By^�rӅ���0�0>X|�~q9�ǲ}s\(�=�o��L	G���݂o��H�/��sV��1jb�A���A�^Ά}�H��L�k�W�`�yQÿ��0���+s����D�%��gӔ��d|9���5Z�LEDSMˏE�+m��%}��ml�����Y⡎�̦��y0��d�|�v �#,�Jn�Z��J*��טF޻��@���E7x�f��1?�cۯ�F�Iʏ\@�6]{�]����rl�I��Lf������D%�g��+�aM%v�tk�X@A���e>���}]�׽~!(����;Ɏ�ތCKɋ4i�gC�F��%Sf�w�S18Ŵ�"f�M�x��8�!o|zQ�d{� ��'^�N?���R�h	�M����F_��|+v�|cC��,ܦk ���+oA��t�?u�^�����I~砫�k)dY�X���k�����F�vz-��qh�Q�'��I�t��,P