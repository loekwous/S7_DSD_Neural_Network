��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�l�(���q�a��8`K�nz�w�V��� P�����"��l��p��2����}�iH��i�k��4'�����C�H-�%����c����ݮ�ƒ/L�o ��RD\���m#Ө���������tw��NA5b�7���ßS����2�+�X~듮K> �1p��M���%���|�8)�"���*q����E�x�-k��A��#����a 0�Ԗ~0Ghg�`,�i|v`����b���I���g �2|���KϦ�}U�+��t�qYBy"R�>D���tx܂�O3(�C�*U%f�[i��V�o���W�R�ѽ�	��Ǹ�L�8hG�]Ii��o�hk=t��zkC\V�P�0�{{M�^<	E�	��!G�I��E��/2T
�qd��HלgҚ������W�o/?Ґ���J|9�4��(:�zX	f���M_���j�)F���|�M+M+�D�j�eB=GF#�`FSF7�M��լ.|v��Ub��r[>?x��IOʕb�����5��X )�^k���q�����'̄�ThC|����Z�F)PjO�X�$4�G$sH~�u�c�p�������}y\V���Ծ!s�ċ��e7�p3)�c���H�V�,�+s����v��1$R�g���x��3	����tD���3E�[wI�P�t���5���#�8*`x�����=�m��e�)�B�gB�S\6��m��'<��#���bta2��[�9n gilZsk���8�S:SE��$P'j�������wM�X��]B�o[����j;^�&*�h��Hh��ł2=�#y����W�y�ʷ�Wd�7X�؋�KD�(gKJ�X�RS��{I��A�͏ЯoR���
�כa�p��G#nt{=���A	{b����m�p�^c=���Na�,�B��D��"��$��;���9y~4����nLܦT�G��'cُ6��8V�{������/3��x�۪���rZF�Fh?D��
U�I �Zܰ�.�A�g\��r���Q++�>�756GO��«�}�Д�����"�s<q��VU�j~���Ba��ZU�����c�e֎�C8s#K[eEc�1c��A;!x4)N,B�E`&Ԍj�f�nS�2��%�Ÿ�~�lk��;�,F�h	�� ��χy���I���7a�D�/e�J�y�ѥ�>��܉|ڌ�y$2ߕ<|���U�y�ra����~l�A��L���\iW;���y�)��tȸb�*έ�Xそb���K�y���NHH�>����TN����eե0�`��Ӵ��BD����D� (KJ�� �C5#b�_T��o�,���z�q�����zZ� U�EH>	m���2�7[U���`Y>�R�$�U^��wk�f�r�-*�L�gr�F��֌Q�i|~|�?���o�����*/qzb+u'+�����V���2+~��f5��6zs6�@���j��hAb݅)E:��Hv���K��Tnei�Z}Ë菒��t�,q��1
��/�ŻD\���5�L w��ׁI�k�1�yak�g!�����JYד����!cb�֢O�e���M��=�!`c��F�A��Sl��稗�����)�����8���)f��W6��rO�R��2첝k.����r�X���K��24狗;�TNqPe�� qM&��2�V�Q�|�ȷ���H�ɶ�p}���>3:4���;�	.�t7��vq���PM�i1p�XȐ� ,A�:���[�O��t������a/ֿ;d�2_G�C��o�?g�-~�9.Q��� ��u�Ups5zZ�f]w~�h��ܪ��8?�K&y-�M̄F�� K��<��t?=�͆3nr[pM����No��)�I��s����K���M�x�=��Bk���� ;	�V"� �R��vnC�(XuƋ�Ǔ+��eykV�3X��	�7Q��nM��	���v�,5��������'�d��ϼ�1+�X�1���,�޳P�3��p�呁��i�;��:�ٱ��~�knQ1�J�`d����S���~��oT:eSṣ�UM|͠�e����;t�׉#�� �,D���,��t�0���_]��1KFd4V/��R%n?�c�带6�`cެ�b��p��� B�&xuUF�y�PjR�F���ͪͳހ�����pJ� �sW������%��k&�׌5�/T����=,7Z�/�B���}�3��W|�Se\�	pE-B�4�E�+��c�E��m\�'�Fl�p�\$;�1mdp�}�ɹ�H�_���х�t�Z����(_0� d�Z�]܄�o��S��G�Nޒ2<�4�/����?��?F����wǔ;A����,��OIU�wږ��Z�x6�vο������qdq:��+�8��U�����(��D�����P@y\��L���E���T�ۨ�>l�g�e�FR ��Ҙ/6��n�sB3��W�)`x��6m]IPW��8����m=E�HD�|�iqA�Ǭ��N&U��I�ݘ��̌5�Jj��VN��|fI��q���S�g+RJ��)���U�줅�E4V ���f�{���εQPXe�1���f�/%�-����C胅��M��ٟ��t�vW"|���D=%��Kڰ�ߴ�_-���=�M�<�C�0�K��,X��Fg�մE.���a�H���!ū0���������~ �U����-*=Vt��V�$���R=|�k�F�
��
�� ����%�x@-P=d�'���nO�l켐޹�wS}-ĖK~C�i��{}#E�\�U��4��U��{GD�Y���[u�a���
m-�q���睝�qMX$o��{�"\:ӒwK�T���LJ3Ҳ��{���jX_a�p&~�9�R��e���@�E҅����Z4�	X�iT1j�j��]+q6�\���.`�.	�L�
�f��y�V6#PS'��Cmaf����A�����r�;��i��B]���,)D	��JMǰ"����*DѴlH; �Z�A�'���s����W!j�Z;��J�l�M��zqk����!1'��K{p1�c�h=�SS:Q'l�4X�Ҍl�8����A�O]�*.�%Z��[�<g����FD�1N���S�������B�a[.j�G�Rb��Rh�)�k����4���4�� 8[\�"��#Nz@|~��5��Oz��Oi��U!4��N�dKg~���#9ɻ�۲���B�l��{y��fP�f� ��o��s�c���1�J�%M/k�p%i�r����qN4�H'��T11`�I�wE��t<?y���K�2�s�Փ������H��Բ���;�&�v-�0��'7���>���^=��Sa�2쯬���0�[����k������F?�<�I|8�$���dBmlCE0�4ؗ��B`G g��0�����A�UJ���m]������=� ��ڵ'ݺ�vݘ�x>n;x�r��t6��0@	�������n,��W�Ś��Jp�"�L���g%h�����4����M ��X!�P�o�}
+ޛ�t��kg�.��t�s�ۘ����/)�J�0�9+�d�,V�/��"�bL5A�j�g.����y�tۊ��D_/�I�m�!��\;���o	�j�o�������+�@%#!�-/slR	5�n����;���7�zSE���|(�b�� �i>��#���6�CC{M��m��v&�(wpJX��TJ{$�e����`r5ZɈ��]�"����Du�m��A�n0o��Lv+�؎0�YEq(I|�w?�����p7�������k^�}I�B���pW���R��t���V--
iRF�B���A����vV�s���aB��6����H����L��G%�Qyr M$�5Q�r��+���Z�����Y~C�߼s"�C���Փ���'�|�m#d��I!��+&�-�@�h&�>M>���I��_m.�h�V�<I��m��^���d-�������.z.T&���/�6~�����NC�>�qwJ.70(��d�ܱ0B��Dkj~�w
������u�N�s��u����Q0Jq��e��~#a�"�i�H�~!�-%�R�2�;b��f'�<�\/gy=�\�TEߗy�got�"`�~�p!�?=I���;#���o�hJ�P�y�$@�p����2���ޙ�3�sjw��ɵ^�t��,���d��3���4�.��W����!2H�y�X��{��į�F�]�>����Q��p,�	�c���YGEF����;�:8��FQ���d�LSz�y�m�z %
��\�v #r�B�6a�RY���A�d�Y��;�*3�������$c��@:��>��l����퉛M�^K��H�S�05"�ܵkɈ���2�l�l�^�//��n����c�;�+�}��D�G�N7�BX�Ϝ�W�.\[=ڎ�o��zu0�F(ߤ�! �~����CZ�U"�䧭?Ɋ�X�HM��I��y���_ƴ�����u��8�~J���ѢJO;�ui8�P�S��`��B�*�G\�h�(�@C�����-r#JD�l���-���J�܈�o6qbmҪ��y��0z���u��a�k�b'��<��!�.���s'2�#� �ngc���fj�����X����5��J��ܜ@�-�IX��� (��Z��1H>-	$�/Y��
^�~�$,�	O󡄫�n�(����Jqp4}��g������a�b��6�����ғx��̞��oD$p�ʋ ֝�����ù��b��A|?�D4�����[6������2L�=9X�V�]��i��"�TϠ��L�����W֡��(X5=s���q_��fU5��v^��a����}|±'�}A�H�^����C���Mߥp%��Η�t�;�أ�(�㊢� �\6A���]�n+�rq���h0��0`�J��~GV��.��`v)�9���)\;�0�gBABŞ�Ĩ��Y�cD	R�d�?'�|'��á�a0!1�͍X�rP��y��D̇���K�I�P���}���Nl1E=�''|���Eh�B�gN�3[�֒����K>KӶ�����Α�g� ��D��y��a�������ܴn���g�v}����֏�6���av}�;d�/�%9ސ�6
����DH7��$�3y��d��!+`zu=�"�X�Q�a�L��>�A�ܝ��U���}��.8���h��B�R�;.Yk�ª���G|alG�j��QXm}�m���j>>֌����2/?��21���P+�����ZB�%[��4�)�(y�ШK��a��A۷ߖ]Ԃ�<��������'+?#�r($?��{�H-� 2���G
YLf5���~ ��J�q��V�trƤ�È��Br�~��:�znR����D��j.;\V�W�_rAœ/w,�s*��|M��J��g�\���b��x�w6;�tDcRY�~@$����,W��s�7Yv/X*����N����p�����[]<S	������M�u�����X� 	��SO/�yH/��޻���&L�MQ6Xn�՛����h�zT��S�xҬ����Q2d�<<Z;A��x�^,:(K�I1x�\�A��)��P�*O��jkx䭟��i'�CQ�D����?�w�_�s���1���W�n"�9J�,��x������%#���cy>㱾<_��lA�[ �_P\D�;87���*(u|�����k�9oI�C�[,�L`ÖmZ�)R��;������+%���*��}/�0NW���X�7*�MIM
3�j��1d���ȀY�0S_����Ƒ� [����:�*�5�E;fgq��,�@ʍ���y*Un���AK>����y��%ҟ��N�
qk7�jf��\4.z	%)��� ��e��E�����9�(PZb��S�0��錘\����ƭǎ��X)Ug-V�.g���MN,�,��^4�|l�,��n���,��K,��Η� S�/�;DJ_Hޔ��a5���Ҹ=�	=}fs} ��l��6��/%_:/���3�7
�@�B�C�i����,+b�2őV��=�?�K�?%�1=��Q\(�9�@��$�$�[���9���_����|�j���q�<�v����*;�~������2�5�wp��z�x/��'��>E��)�Û1�8�����a�w����*��Ys���;!�Nx��{�ڈ��:�*D}J�w�\f2%[�:�+_�H$�R<���,�+�[n��N�qb}U]a��U5G5�pX�`2t-|{9��g��g]��O��m�|�u����`�ZA���t؜��e��[�BE���#J�yk-3�i��� �2g,�B:��p�R'��%�\Т-7Nl�wY�ƌ8�+�5.>�*7��>��}���=�`��U�m���]��R0K��^�pm�ђh���/L���b �b
���D`���l�X$no& j�ܮ^+b5�%Dd<>=��%�Ӛi�t�0�;'��"C^� ����Z�w�������b%������2�MJ$QyRZ�q��@D��"J�P'�v�j���T\A�PW�<�7�D���\ɩ� Ry��4/�Ux(x�.��	28��)�.9�X�L��V�Tt 6���`x�?��dp�g=J�����X4�i��0�3��;�V������h��*�0�-��q�)�c��"$��ڋ�.{��[��d����!��q�����b784� *�I_��)i�*�����m��0��=��WAw-;�߷�^[i1+��n<�n��� ���,S���=%�*�V��VX.�N�9�pnf���U��H��GM�2��#����<�Z�61n�Kq��.��=w����*�U1�Q;D��9R@Q̾�m^�&�y�⯯����K�dA�Pǁ(ڄ�0���
�����Ӟ�3)_�*�^T:��[�Q�N��{�#�.B��o��1�z���s#�D�`)R=D�{�E�s��6�`컎�%�Y����~L��<DD�rwZ��D�O�̎-�> ��3Н�	�0�u�	e$�bkJ�E�M���HE?F��Cd�P�>�3�=�X�8K<i����J:����M�t�=�!ܶƒ�A ��.��w��������'�u�P|��7��Ym��PS�R1��	��X���H���jd2�u�s6����qx��z�.��M�U���=R��D�R�Y��$��)��/���9-��O$������قZ���Ҫ�>���6����m�h�iC���������dQ�Ta�����y� 0"4��:'�{��r#'�t��4^�I���/ի��#e!Tټ�̫�˴X���s�I�t���m�M[�:\cE����El�H׊���)�E�i�
A_�oLVG�[#k�j���4��dS�+_7�̊���Q$n���Lq���!�B��h}�)�YGR�YM���MO�k'5�)I���t�q=�=�]��_��NV4�`h`�%HG�i���E��*����~��(�jG9�:��������H��Q`���7�5��e�Фpf�x~��w���h������B� ����і��Tsf��"�K�I�tB�����Ut�}���n�bU�ë
�a��#��o�vj9r2a�f��X�&3#�V�P�
mT����w�2ӄBD�̑F�_�r�袩�7_x�w���/�צ��7��,��dҗ��7|�J�H���T��*3O�X�L�1��I�}r����c0#����9K��4V�!5�x7�]±Z'�fq��Y��x��4ګ�����y�}��W�U�Ϭ��xV��[A�����0�"j�����&�O3@��tyày��ߘ
8g�߳�4F�<��V@�� DS���cL؜b�1~�!��!N���E�����j�
ϣ:�� ?���F�@��;�׋���^��7׶"��N��ȝ�oa"T��X��������߱�LBe �R��G��.y�`^��)n��`�_� �#:6���q5�l�#���*�7%t��E@�|Ւ�y>���Ռٜ9V�}���ȵD�-GJȍ�ˊ�<`���'`L��#�c��+�Dm�'~,W�z
ūe��~v>?��;���'�lW����|�Fg���H]�f�b�vQ��w	i�s�oz��K�z�ķ�IX,T�����=~��}�u(���%!ۆe�� �
[^F�3���_5RlD�%]l|��@+�i��dp��4�k3t�ag>;I�S0P�$%Rf���S�:�׻�]T{�"���Τ��� �~My�छ�XTB�l�Y�
/�&,��ܬ�y�c�q�1�+�R�׍//Q-W�������)z�4���z /"y;�t^�r��Y�C����S#�X��r
���W?������Y!8��jWo��������I��ra�V(=l�`b��h��'�B%Vif�T��e�P�xYغ�4dH[���6
�w�e=�:���7��93y��3a%?Yq(�/(Ĳ�%9'.*&2��6��Єm��6�d�d	���2`D���~-�D��6K-���V�uj���Pu�7�̝^��]�n�]**r\���,�H�r/v�$����FG�/}`��!5���ƺ�¨�qxf��$~R�/?!�6� ��ܛBz�e�s!N�Rd��^30�O�L6wZV�f���_����±Ȑ�<�?}�ҍ����W������z�f�M��I�V�.ċJC?�MI�q�f�I�}���v{0�����GF��oћ��A&~�o7��ܥ*���L]r����� ��N2d�÷6-�br���}�'�F_�d K�E���'����-o������7\�~��f1p�]t��#�ֹ�E`tө ~IL��;����%Q)���f���o�����H���5H�4�%�kX���b7��L����D�B�B�)�0�=_�@Yh>��4�i;��S};��_:e�π���m�^�h�V�t����q�ǋ�W��3�7A���y�6{9�����cL'�˾�"����-i���6ѭ�;�խ"���8hS���Τ��ա%������=E3ZpټA�5�4R׃k^�̮u�AF`�h�;�eE��$t.��7-m����V0�r���1r����j�?��2�
ڊ]���`�yQs�l����ݽP���y�i�Ӕ�5����m(.<�%H����)���m`@��]�Ѻĭ�L+����Q9N�-g���:���dd�黊�=���vs]J����\��Խ�]$��(��L	��9�A�������0����>�B*f@�0�s��
��]ٗU�����B��#�[NǾ2I��BP��+�!����(��أ�껼\��|��U�f�ճO��*O[��s(Ă���<׍�f(�vXX��=QD�5�2]�	�lO��R{
�t��.���~�&��SJ� ��2	��w�yC<n3�T^��.�#>μ��ؼh�>���}__C%+(��{#�w�ޓ	����V�ZT�r��'g�z��i[z|ЇieO�ᄒ�z�<	��_9!NYK�U��/]ic��&�����1F*	nF/�Y5��1�;Eꞗ�ң��Y޴�����Ǵ�1�-���B�w�ȟ�Z���Ek����ߊ\a�<��-1�`�9�W����Sږ$wL�$��s�q�AٱX01S(.���T��w����;1mwX3DQb7�}�a�/=��� ���.�W�����b4ʦ��#ː�k�z��$���'�,��(oӕ��f���!�n�U�'��{��9M
6&Lj����� e8��#ev��[X{�+��*�D�mX���Cp�Y!����mK��>�ۭ�^G5t�,s����:M�{m����P*�!;\���A{��;O��v����y1�-�Qu�r�h�D����>k~��e��f�j��A6�C}�i��S\���*�.E�@l��^J���v|3�a���t��$Q�^���rm���PI��M}�eÞf%@���*�o�݀�-�@���L̇j!�dʤ-dV��y��B�T��Kg}���`��',������֟�pn"��鳻eRN�t7��T���l��v�� $��RD�s��F��X����YO9�Wf��)c�~#�O*���M�E�U�Z��7�4,きG�>-�[���.�`@�� �0�{�X���q�G����R�S
�[YP? �Z�!����0ɫ�խG�Pn:�ɬlv�ç�o�o�h�)G0B0N-خ�y����Gs�Yݧ��~�i���^$O�:h�LW�A��nV�(��G���V��BX޴K2ȡ��Sqx)+ì���*'bO����Փv-�0&���;�G���/�m�\�G��V{�V��b:C�֬7̝��b�/D�h��(�k1B�v��7�d�� 0kc�����T
�M2��h�
i��ѓ�!J�����$�}$�v�\�eM�n����@���S���$����ٸ�W��kx�4ī��@��^'P*	�Y�t���؂��O��(��9����Ъ�%\����Ȗ&�� ��4"���X����)q��#��ؒ����s,C�a�s[�*�3ٲB�E��K��O������Ϻ��"86���c-S�2� 0��~�Eِ� o��H�c�|K\��Z���]d�����J�
�6J[F��󒦧λk���а�n�Fa��c�g�?��J��!��j���)v�'yt����8V�xq|�n��s5��^�w?��K�{gj�H�J^�k�����̶�K�}dn1��v��N� ��z�0���=Ɓҥ���f����'	��� ��س�[<h�1@䛜|��`&\ݴ���`���ռ�����[o'R���F�{�61�{t0�_�M:I�b9�ּ!9id.�h�UK6 ����� C/��7��#v ut��N���<g��?h{˷�屒l��jr/���t��ZQv:b���p��B�V굍Ja�3�Z�ć0����C#J<Eb��J[��t��sJz��r���_�E���&��eh�z�I�M>T0ʙooWi.�a�����>��AzJN,0(�0�_�Ќ���N�����J�����p0�S�KP^0�m�ί��oTM��𧕷�2\z�|
Ҡ�eU�l��'>q�^�I�B�F�?��J�~Yy�G�/jp��Z�-4g���,������<Ը�b	�ܔT�a����"h���g��oԩ��uHb�9-�ƿ��w�%�H,+�u��\����p/a,���H06]���3K�����M�҄\R#�y�_��n�?�^��VƳG����~y)���SK"m�:qY@Êm}WV�5FA�:�j�`������^4葼��2��N�[A��}��T쭦�*$1Y;�(����Z��t�L'�c#h)�۽���Ç����YEo�f�)͟���د�ZNfߥG��E[D� ����g���B��ǃ��,,ѮKF@�jԟg��G~��B��Ge��wfD���bRJg�.�0�.��ԊH�B��Q/����.C�e�ƪ?"��wu��<���+�t���Aİ��l���G�ZԹ���u�sU=2�ͷ��'��/�+�MO�'Ly�_}E��j���J�P��w��J��v.q���T{8�o����U���)k��-�1��V�!�X��V�#Ɵ^pv�C�BpD��h*�s�O�ᖃ�����Y#Ş$�3]��^���
�C��*��c�	�n4RU.y6�M�g �j��U'�-N�4��������iTF�jw��T*����V	��6vM����.�(� IW�yS����K��43X���ݴ#��k�I[�J��0��U;f%��5G�>����ѳc-���Z;ι��'��Q�ʶ�R�nGܝ3�>��yS2E$祌l��zD�����L-B=Q��U��S���O.�n��HO�Pd��|�WWh�b[?</�nN#A�l%1�I�!�w�7f�P��Z��d������"fP���j�R�DiWP	"ԧI�`��#>Si\`�9�����"��)�
~���ho[+��YZ��Î(��������_k�S�OL�1�^�dH��?�Y?�D�^��%�M>���������"J2=3O͹-VH�F�.ϛ��:��A�\�-��?V�����&@G�vQo�ݽN�q{�l����jVP~��&D�J�,��3T�Y�B�ÁK��Eم	�J|�L��k1t���S�T���0��pN	��d���\��%���$��|�nz�e�e�d0�Q�xc��7D�6��\��c(�`�+�S��"�ֱ�t�1g�>.���,��x����T���y��O/�S咅��	�)��?!�뻡Jx���Ds2���)Y��)Ƃ�yFb=�"��ru3%�g�8�e�yS�6xQ,�� ��}-o�D����n�e ��Z��(rJ
�6�s��Q�h�
͋���S+�����y�$҅_�j�Vx&J��|K#b��E�Nq&�����@@���c���t��K1t�VM���4�T�#�S}G��� CS_����5MJ(�W4ꮇ3�K�ň.���Ȁq����i����|�IV�~ǟ�ф3��X�[�xg�f����7���K�?>��=LRK�j��^�6�o�~�0=zQ��|1����>�*���6�~o��T_^z��V!�	��A�fD�w=	�����J�h�P�i)ni"�ۢ�$��:hsk"Л'�V&eI���~5�m>�q3<���c�F�`�6  ��a�fcJ%i�I��>fvz�-A���!��W�N��Å<�"z�yx����_P"-_(��ĥ{�2�x�)�y�� G�oL(�|[�D�RD�cM{%qG2kR�s~;�Hρ�Rޮ�a�v�t']��QWC˜��6I�1¬E�c�e��154]͹��A�������[gr��'�wOm��6/�sX�����p�X����4z^��a"㜱������}\���1;ڏ���I��M��͘���2J���� �K��Giלq�u�R���<T��j�87���/m!|-V"�f��/�z��Woc��l�`��2l�	*f�v�ݓT�:�]�PS��r�ϒm�k(��a�t�m�fZ��y�� �\q��v�+�'b�R��Su����^��q���xu�D	�:6!�N�H����9��6B *�a�ff�+d�Ǹo?�R��*1�M!=�x���j/EZ`�e62�9tF��0Gˉ���s8;�	$CB�d��e�LL��[�.t��w?�sQ�3��6����N)OE�6n��N�z_��`琎J؉|h�L]�U��*a�~0�m)�xm$B׼��tT��4Ñ�J���nJ�N��N�U��.v�b	�f����%�C���KH-�< C�*�\V����DҪ0N���LW����rŜ�?��kEh�o�gx�����	�2�
��g5���m�jb�����,��ÿ�M�0��'�1��D����:���y-#���L[s'r5B��W�x�wכ�����/x��[�5�Ce�P.JdCzWb_�l�3A�����qKTPyE�߻$�Q�"���$���"��� F@�2�-#�j��}M�.A�+�_������0?m������|��0�r���:�>d�~��^��'u��Ԭtve��.Ծ�F����*#\�r��Rwp���c�|��^�|d�W þH�z�F��N,H�e�$F�Ř��P��A3S�Ƃ~z}�)9�jB���z���r�ED1���Ej1crz��"�����"�գ#7�ʱ)Q����l��3���g����q��}�AΦI�3��
�5S��H��й�[���"/�X1�.9�8�t?��[@ăާaa����D�E���h�О�!����4^�6��N�e+.�Uzv|jAzW. �b�YG�c�h�_Qi�^~�;^�>��3^���x3ya>I�[I���$�
m�xJ#ƽeR��O��So7f�G=ϫ^�bSe�{���.��H$��w���~f��Y�YP��حX��"l��x�5���7���>�: �"��LΤiKoܙ�'�͓�ßz(��	���EȨ@-�e�;�
}
��oC�����Qt����c����#���Z�Mପ��xVs�>���}�C��)��
u���˻L��$�
�@��=:����g-����˅r-y�t8�EA���� WU;����P�Ψ�����ɧ7�|�y$�]�E~�*x~�Π1�c��rLc
p��c��K:IHz9���a
wυ*�n@��tU#=�Ǝ�<SM���H�o|���Z�������s�{ǲ8�������s�o�6��mCj�߽\��6����
xQ9~1�� �d7JC?G� .�=UZ��k:��⦿������pX�"��+��$w'M�I��]����,ķ/
2*9�
�7�A��hS��G�.�:J�7_		�ܟw�h&�Pf���r%�%���v�q�]�.������	^��ۜ�W�l�Y��l��I`mv[ �����Ľ�}������X�8#���=*�S�����勓T�w(*�T�j=�/4dlY��l	�Xz�T�?���F
T6�r�
��O�1;�y���Q�%�n�z�����hg'��?�m�>:K+�8& X�U�b��ܦ1p�����6�@U�kcN~r\I����Z�}M��D��F	<T�٧[-��#�bײ�K�m���RP���%}���a����W�L�5𝤢,j������>��.�����ˍOB)���ieH���	L���*�:D_��h�$v���x��A$o���mx��AGDؖ�ᤔ�-S�u���+����/n��5�n�Li,E���G!����5L��^B1x���om<������'ũdP@�Wd���=��n-�����Xu�U���]!kА�Mvj︗����2�_�����8|x���P=�ޘŖ�BODCPÁ��j�ip��i�_h���]�ǁ�\���k�A�9��hE!��IⶌA;4}i��J�ψ.K�wy�-�X���?C��ƴ#�ʸ����W��-�t��ul��O�vۨ�LaU6/tJ�"u���[ܡt�!}�L{���������������\{?4ZB~�v9[�y~1T`I5��S,�q���+��)X�֐�5��~]*Z�2A��<RR���� ��M�H��q�y=*�ŋM#��Y\�lDh����pS�yoc� �+�X�SzX�	�s�@��'�fξ�'���A̠=	�$���.�_a�hХ�
dv�Z��-��~��e���O;��;r�v�
<]�È)ܨm����n��V/��K�AT�� ~�A%��0�\`$��"���޿�L#�.�dI�b�HfK��N��}��})N�,��'�+aH@x��aN.��<����=�އy��9�c��f*]<��h�A��)�o
>�@�\�`U�	,���m�FT��.*ǓM�C��(��C�ix��Xb�EV/��A�z��A�@�~�zʳ� Ʋ��y���3oQK�C��fN}vW*�����6�P,)u����vx_�Ꟶ/��@�.���HU�;b�F=��]c�@�F��� '�T��f����>mC,F�g�aR��H���q��د6@Uk��~�1÷7^iZVD���ZZ
B'89�d�O���hUfsz6��}���yF�|�|d��6H0�A	S�3P鞯��t�4�gu��!}�Y3;qh[���E��僕�s1ض
�O��B�]R���x�f�X�;"�Rý�T�	YV��� r{�K�5��=��Uu,+�
!�⫌�ko���v���h�2�0Sj�y��'�]v���m�����D��S���5���xm�.E�������9���'>	��F�-֘�H[�N�Uç?��k���g`S�{�7�<��~柒w~r�:�� ��^�]gB婴���:t~�|-�����c-��h��z�l�.1���#�v+�嶐�S�D����⇱�F"�Ǉ��D����TK�v��P\&�'f��jަT��=w	���s�z����oqڷ&_�Z��]��G�kڐ:NwnAx�G��|��5�?����LV2�Z$�z��Y��wu��`e�F��j7Z𫛺��`�
u^��3�4o�[��!Xj�@<����kԃ���'r�?X{�&���YS�<�D��UfZ���o&�o_�Ó���%%=2��-)*�˚k�V��~�k��#�<I���p��P�7S�}3����	2�>�g�\��ɶ�IIz`*}�khʣ���{d��\�ь~7fiH������*bWȱ~YG���j��9/[�.eI�7���u�2��^�H�i�l�3�����iL(����C�@�F�:.��M;;_�}I�ݫ�u�A)��aX9ÔW+1W�(����MN�|Œ.��[���M8�i���ܧt���@_ԉ]�|�BM���;N9��
-���	h*G�ԕx��pվ�U�xX�\���H<�n@�Q�ps�n<�Bdw��ۘI-�A�E�n�7l���wS����[r3�[����$�K�>��GGs�DƜ�fHnm���M��7^���<��=2b��tU�[�Ai@o�xJ���%1ܔ^HA�݊d��+�z�?�5P~� �(�c��6٘}�N%"�6U�������}�����?婳 �C�v���g�I6/�o.�����%�ߛ��y�|i�/����go�� H���18��q(�5p����FӸ���f�>��@�۵8kY��"��N��y����cq4���5O�G���4
��GkF��<{׋jԿ��7��/m �R	��n�\�4���C�'�$�H�J����cJ��qD���|����]��%�t��:p
i���	����A��	Ǳ�������X�1��F�����H5�!KO�����q�;wT���)�ΓX��D�a<
1��>n�]]�H���_X��&\�?7|N>E	�l�c��en����
�WLZ��W��ǐ�ԁ�#��G�c!��{j�<b�
M9%����j+�G&FF�I��W��m+�I�Ɏs�u\:c��8B�R��i�ph1p��W;���%��:~�T��I����`����J�Ɣ�,�{�8�n+�{N�����=r�K)k-ވN�:��=�T����k=+p�
r��G�S�#47�}l B_�+.�!\%��`FS�a4�h����hR�����݌�Bۃ�#ZfU9c3�U� �W�������! ���Ťo�y39�J8��*C�G"��;nʊX၇���C���0]E/�ϻC�#V|=�@H�m(��ˬpl(��!O�'��j�y�gz-ؼcbi�81��5�c��8���&�m]y�8�������<)�D[y7Ϩ;�T�8K3ƌ�|;v`*.L �(�W��
 B� f\���wV��d)�v��~BV�O�5��;����r��f�߹f��YZ9{D�Md���[�)���+�fݏ�
K�y�c�A��x�o/�C|�c�K���mfRAjA���~�`Y�%o~��ϲ��1Ut`ޖ��Q�Gs�z����R�Us�Cb@�姛P�Ii�`<�������i���v�;��pp6�I0�]����)w��`2P��Rc�-���'��Wr�jwjUF� �U��TuX����g�tan0w_��4XX3��V�2 fT����)�֋YwÃh=��3�(����I��brnn�[\Y�ۅ���'u�'�N1 �P[2��:R�5KrP���s/�����q�r«`��53�k*Q�;���~صE���i����95)D������&8$c-���(Z+t��U�[�xD'ǩ�p�Fv����f,�ܸ����)3i���tlH�����C�!���r'��~NA�C}oD���R}��0�V���;D�u��?4\�M`�QZt���O����(�b7ǆ�Gu�GOΆ9��}�X��Y"q�P��k�&�W�ذ�MViB�o�۝�p�8Ճ,�
����G3c�)4�w]�p�Y 8�?&��g�����8��*tw&�Βېګ���o��3���՝���i����"����m/��0:a�eg��i_9�{��	�7Eg����8����H��xo�O�����2��=�ٰs6�A�
��1�>���X�՝��4�,��_-,
�pE��NƘ�g�GR��U��V�I�]RXPh\�H�i+_[��p�����\u7	y�R��Q-Sb_{��v����6Gֆ��`4�J3��1'�<�jG���� |�q�w=�F	*���9��v��S��x8X
��!�:�#���a��)�j�eWc_��Z)��g��Iu����c݀(a'%�,^4j|	F:����#�Q	�D"[�NVX�_�@�a��Tm����W�{��p���]��Pz�#�.�Zy�3� �YŹ�� h���۶9��J����@�EY? [S� G��kMO\}j�p�+�yܿe������M,f��q���ăW����������P'_7cN�0]V��b1M���*Z�-�
Z�N����_��q7�\���Y�P�_5�F�9��O�#����|՟�B����U�;���騶S2�����X��]vX�('˕��x�h��-�42<H����_���
ǃ:��%cIy'�J�CO'����z�i� z��
a:	�T�rԸLɣ��
��C!+��Y�:���)%8�%��r���!��/���o"Y����
���K��g00�M��Rˉ���.r�Lȗ����߂��@����2Û����A�Q�1xN�O/��ъ8z
ݞ�֙�Z�ܠ��R��U�o����ʱ�+�|B������1��u*=u��*���K�����g�e����w!�C�N(��$�z~�PHw� E��	�}�}�����V�-�&}ڣ�DAgF��կv�]�Q�[J�j��\���E��
˫���=�}I�}���KpNm�=U{��{�-u���C����h	���9�8�3Nߊ�O`�<
��8�
����`5��Q�^���x�8�!�q�'��N�S�
酒̵vЬ��e�e���F׾�%"x�.��P�4�xol��[��>�h��$~t���c�,ج�0]�g���wԁ$y��t�O��������<=3tC>��B�Ƌ2���G�=�'��q��ep_Q���P�,-Sʨ��^���T(����|�����!�b2-<�9m�u9> ԅ~0CQ�c_��"29!!u��E���±*��������u ~���^����nG�؀������F��1휃K`{Ff�D߿�����1s̪��]7M@��)�����R[�)��vf�#�Sp=*Ƴ���r9gDE�Ud���1@s/�K�6J����5��G.1+l�����b�t�Vh�v�o�#kĲ	������xtdx�w~��ObF�؏�wf���G��ԼF���^}Q�� ���!�v0C'a�>��t�|͛M���+�MiyT��|�mֹ �t4�:��(&Bٞ?���N"�u�3j^`Ǽ�5;1�}�i�p��z_��Ͽh�tv���/�.�f�ܛ��3
s��G��=��k)`�A�B�AۂGqp���P��:��(�C�(��㯑ȿ��di��e�`�X�E�����$��Ө`?����L�d��D�'�>����m�]�NG��ԍ�àc�k�7$�|!q�{&U�⠣���[��9��V��U�;��'�o�>�$�J�|	Xy�ݎ1�c��šI�.��n8�!7S9�a��ƶL]Ğ��q�KwIp�nbj�(�� N���srn������PT�,1����ݳ���]�zR�dp�-IZ�}����<���!_�g؆
���%զ-a31˵������\��[�=-��;�c�����wf2+[����r��wHi��k2����v܌ \�5�/��FĜ�� ���P�J��h�M��)�&�h&��D���>��xZ5j��Q�z��,"�����Ťk���q�ޘ%����4������(��5���	V�g�0�A�O�G�e��r1�0��s�����}�������p�-'M�[RA�f��#nӖJX:k����[?]2�������$����;u�vݶӫN� ҃5r�*_�	�1��QM~������Ћ8N��g�Qq@�3i�PA9�� ���rP~���i�U�(v
��Y��C�^��w��15�>��&� �[~AՒ�#3zW��QBH��,a�g� �~���7��ٶ�sݸ�R,z�g+ ��T\\޼�~�w�l����cs0P�!�K�+�{oi�x��Ǐd�{�"��Զ�����4�Ӵ=,	�W��l�~?I��n ��(���Y �±ץ��BZ�ű��Q������R%+ĝ�I\V��b�[�bI$]�Ud��վ��􃠇8�Z��G{� "�RD� �������I��>W16�m�M�8���ˈ�����J�ߖ�����S��o�����ᇛ�����X��z��i8�a���%�
��{2ꭉʾڗ'������+���G����ŅH��u���#D���#(�^�L�4}-���`���чӷY� V��O��RW����<���U'fw;�,�<�@�lڛY�1U��?e��lРL"(��|�6@j�,#zo�nN]Cz/�·+��#9��tA�<����<[�P�[�*�ד��ڛ�۲�����o͜JzP��=1h�k� ��6G;�c��� �Ar�m��?H�M֟��N�VDrDWTK�.��o�6��h�"��[��xV$�h�����X,\��I�ٰ�O&_��#�b�4���B{���7��)$Rd�]>��l�f��29�!�efOhE�DUW �)h&����-��}j����"�(�UR�|�׶�h�h�iq�^P�6w^�Y9"�ڒ���l�	9T� h�L��IPW� Qn��Nȟ^kdv��f���.m�j�X����-�f�9��6�����ڒ0j?�*�y$o.�[�;\+�q��)׸�Fɘ�K=n��[�X��r�|h
u��W����ݜ�6�]�8=q;����p�o���O��O\+��x�2=+;?�¼��?�4���V�$��]�N�r��>X���Ɂ�:�*��T�޸IV.jS�>���f��+��F�%Ǎo��b��G�����$�r�ψD��MKZ�x��}���R��2@Rc�s�@��Ҧ�{�K,�-�ٜA��(�h'������ĺ�e/?JHf��}���#�l�s�eg+�O?��]8��$�=U\j.H�냟�Ah��,N�^S�:#wf��ʌ�8uY�W*ͤ[� M$ardR�r���T���ү�#��ʫ��h>��}�� �g���y����>+� ��@�3��FK'"j�G)97O���dv�N��1���meB)���L��v�а�z����,܊~�#ǡ?b�YQ�����,��;����!��~*�wඁ4C�]��Νʷ�L��\�j}/��?��9�����PME�T�Ooj���	�~~c`��Ke��_�/�Ysp��U8yi�tO[+$5K�����������DQA�Q�yUt��t��\�P6>��n./�Cy��8��Rۙ������lknOD<=sk����5OP��rQtsB=��6��n���}�Ŵ�5An��ڕ� 
�1�\'B�.���T��;�:��u���� ,�Օd���&�B��{m&�.�ԕ`�%5
�yox��*oW̠���{1bּ<C�Q�F��]�~��*�m`��e��͐O�((pm-�]Ky����I^�����_������a�],�����|t��9�?Lu T�؏�M�����n�V2?ۮ��&�3x�u��-��ԝ�)�n|$��S�L��>�h��ϥ�v���ynZ�2�"�`DV���u #�		��uj�n�Yp���3U�����ܛ����L�p��"����3t`��;~s��*R�+}5���Q=��!�7Yy��,�@�캔��W��Wdv	�{d�>n�����>�1�:��%f�#�_v��&^vS����[�c};����ŽW����ƴ]�BQ����G�����`��5��z-��޵P�G��(L���3���-�@Z,�mC]p��7�Z���L�$�t>���	kr�x[#٭�' �xp��#�I����]'�65.�',�䂳'A��v8�v�_�CD�����3������&=0�#��O�_��*Y�KB�۠��4"��T�*,�=�G`q���V�t*^�y�Ά��hf�&�Gu������vrz�i����V���gT�����jz��b-�9�Y� ��]Xc, gS����	-o���?�������JA���i��k�(�33�BX/K�H.�"z����eE���ݺ�Ĩ�ͻ҇�F��r��,dRA����/�L�fgx<D��G� ��`j������A��^$��qlw���x����Ĳ/������1`}b�`^>��i4mcd�r����-�;j�w
y#�U�`�]���|,]��㕓c^1x(�ʳF���&�b?�si�WF�&���3ps�Ɵ��x<�|����q5:7�,v$#C����^J��6?�@fN��K�j�;�|��639{�˖�x-J��L�n�y-�nѸ�B> �ј
��6CX� >G*�{Ľ��uS�&n/����\�;f��?lY�� :�7�Z6`����h�>�����pt%M�h�����W �@�#ln�m�������p*��jĆ�A�ՙ>NaᓒJI�W�|8EN���!(aI�2�*�Y��� K�48�sR��/"���ʥ�Q�И���@ŉ�s�