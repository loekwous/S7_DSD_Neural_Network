��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�l�(���q�a��8`K�nz�w�V��� P�����"��l��p��2����}�iH��i�k��4'�����C�H-�%����c����ݮ�ƒ/L�o ��RD\���m#Ө���������tw��NA5b�7���ßS����2�+�X~듮K> �1p��M���%���|�8)�"���*q����E�x�-k��A��#����a 0�Ԗ~0Ghg�`,�i|v`����b���I���g �2|���KϦ�}U�+��t�qYBy"R�>D���tx܂�O3(�C�*U%f�[i��V�o���W�R�ѽ�	��Ǹ�L�8hG�]Ii��o�hk=t��zkC\V�P�0�{{M�^<	E�	��!G�I��E��/2T
�qd��HלgҚ������W�o/?Ґ���J|9�4��(:�zX	f���M_���j�)F���|�M+M+�D�j�eB=GF#�`FSF7�M��լ.|v��Ub��r[>?x��IOʕb�����5��X )�^k���q�����'̄�ThC|����Z�F)PjO�X�$4�G$sH~�u�c�p�������}y\V���Ծ!s�ċ��e7�p3)�c���H�V�,�+s����v��1$R�g���x��3	����tD���3E�[wI�P�t���5���#�8*`x�����=�m��e�)�B�gB�S\6��m��'<��#���bta2��[�9n gilZsk���8�S:SE��$P'j�������wM�X��]B�o[��O|�TD=T:@�G*�6��B*�>{��
1�(e�t`�k־'�NU؝�"��!Y���泤O���a�:fiE���s��r��Q�,SL��Wr�$�	|��S?���!"�`�6hp��rY�;3t������m��j�����%@�6z������;˧�U���o4z$1K���P@[��;���W$�.	D�K3�p@uF9�yHf9���L��܍��'�dA�\, ߿���&������ [���i�qF1�sd��al��F�n馷�A_�²������=pL�35lu�Ͻ�ڹ:ذ�т"m�Z�^��eb�����/ntY�_�Omx"�֍#*��n��By�V*b��s�n���i	�A�[�\��'����d�3H�>h��Y�lM����&�AC�ҷ�k�^&H;�@t�z��jh��cg��LO#��*؁(4�j=�Gr�
�Vk�H&w���@������6��K��;�6d8�<b1u"���s|���8$XV$,;^����l�2���s��?���M.X\{�C���z��h^�U-�G���t��3�5����_Ԟ�.)9}�i]���4f~�_�ᣙD��&L��t"b�4�C���p��v�� �~��o��U�Y�x�L��*������/����B>d��6�N��B�l�9_E�A�.�ǽf��;a��6��*RA!��l+-����UiP��(�\F��g�+������g������<־� {���{�D�D�C��ӸU6Z^�>_�"��G��*\��OWV�
z�x�í�fh�ʚ��"Y5�o9g
X�1w5YdŘنp��I,gNp�.�o21L�#��=�@Ш�+C��\w�:^�Œx��w.ɤ�ĕ�H��:}nb/2=R4���O�pH��Gns"��fEKu��
cuJ��'��
�&٪]_�p���R�NN+�i�������!{�6|� ��vdI�j����"���j�%`�HW����ea$���K���m��A`:�&������s���C���� ��3*<�U;�p<����qY�1Jd�Dq[	SM��E���#�נ1*o^��M��%�,Y�E�HO��&ֶ��Lc�X��F�r�u���2�r�0�������_�A;�������̐�I==�t�5;�56�U�/��Y�Q��ׅA�#�� ���9jK
���;��?��cjI����ů܉3�P�=h8���t�TNƁ=�v _2D��_cm��蠋�o�2��v9�	$����l,�����-q��~�;�����Ee�a��~0M��g�M���V@�;�������~B2z�V���q$ߜ�!�g ʔ���g~��P��X_n��0-xaUUҾ��i�&�ș��Q/Z'�w�>
��`�@$=fy�S�uhdHՓ���v0��EF��#��LN�ȇ�7�p�OG8�o��w���a���\���������b���*�bFT�G@�w�7�d��ϒ���;y���)�v�Ϯ��,$!�o�~YԚe㡼M�>j)~���=X<�M���������O�ǃE��Y�fK��ɜ��.�.��H�N[`(��8�m3p'��y�H��E�T�j�s�Q ���|�@;Ij�}�)���={F<L
y�\6Ԅ���S|x@4O[e�^{�����ʙ¨���Q�>��b�0��s���J��-8k�&������΍�le�\+�ݒ�1[3�5�vJ�.�gpIu� V�3	���TβLZrH-7�"��[�Œ�$�jVQ6q,�}��w�O��kED���:AOn�Q7ߤ�c|(	�̸��B���y�C�K"�`�dO�'�i�9 ��5F�B��dCK���'|`��������g��I�8)RT}�gL�����v��rfY���O��F��E�q2���ڜ�T����m��f�8�x8WTu'��,4T�$����S��D��w&
���5����>
$��-����T�R:	���_A^��G�_Cs�nNC�Mh�J{�����$r3Nb�����-E���Ax��7�n����5�m��CB`���Y��B"J���4sƸ��	���0oF��4�4�aB���j:Bi���LM�éP�y:��r?8#}K���5��eh�R�a�<�7��"e5�d�<�:�Qg X@�6x|�
˿5
�.�q���1�˙���8j�#]���+�y��5�A�1�;��!I������"r��w?H�D��d�(:����tc�-��}JL{w�ذ,�_��y��u$�؞���s=�eJb�J�K�u�����0��g	S��c�{��ר�=V�Cx���g�V*h6�a5g/y�gS��@�>*0�������p��� �S�C4M��*�ےk��̯��ʎ�c�(�r.�R�{lb��QV85���d^xڰ��느�+hg��QR?�s�
꼑!�1���~C&���3tYK+�g�L�'��4��a�\ Xf���1*�E� g���r�:נ)U�-ɦ*Q��04��\�~+pÆeyJ�i���������3K?����pzt�K/�FYXpHY�W̮IN��>Z^��UW��O��3@1�5�O7N
} S�"��y�*���@����I��ʰ�G'Y��3}s�4D� �q�"���'j�1���s$�궵���uѢ�"ry�\Z��`�Ԓ�F� �v�n����6sȩ*����(�J����O�\�V]�O� ����n�M!F�A@3�@�T$d2+������tH���֎�NQ"0���g�1N�Ze�yÞ�w�$�kzSA����W���������,4���x�`��QL� m�2�p0xQ �A��sj4�?/�
�:����!��	����ἸQ��xonE�4/:�A�#�G��"?wD 7�^J�^N���\�ܭڶ����I���G��"�a R&�L���u��1ӳ[J�	��o�F@��-7/ �� �1I��u LSU�F�Ep��
��=���.�䲜X"^�-B��7��)�ZG���+���6P�R�l������g���H<��E<�+�|rK�[a��z�y08.bܺ("+�\~3GT�I<�(�dN���1퉆�Բ��ow��yr��R����l!�� ��c<���J�d��5������=��3>�D~���y�����V�f(�B8�;o�m������";6�#&�NeT�|�{��Ur�àq�i?��i���ė�95y�3O�H��<X�L-��w.��'ϩ>�A�_l�A`�
=(��4_|^!U�B�`��|��@b/6M�Sg������GI���[��ٲ3��4��*�G�W�R�1n�d�eB�v
G6�-�
!�_�:M�����2��v��҆�G~�b$�9�����PA��j Mn\����,��.�يw��px�,��zZ��2F����k���k'Mp�!#p�h�͓J���5�]>�2cև��DǠE��Uv*��i�U&g= J�|�6��?�,X.�3y�$#�>�-�''�:�&��z��O���{#�s.rDq�����i�T��J�	��C]�O]��k�
�bdj&��^�Npl���k.��X�E�(�q-Y�I�n��ݯ�V�������n~Rs>�x$G}ʘH�����^jB;��h�W-�����v�`�:Y饁�r�1)�G�QR�,�"�U����c�U��cr�y�)�7Cl*!�S��~�]�;&!�;㵰�.������ز��^γ�#�����H����fO	����zM+;�',�}1D|�y$O(N_f?�1���|`1
��J�����{�4z���p 6)�ԝ�,���r���ڻ����=v��bގ��$B��gӔ!;����9�W����I�������96���Jgb����'�-��$��`�
���� ho�z\P�Bi�ᴞ������������)��]j�X5N#B�CV7��܆ R�=Xx���\,��W�i�ïD��*��	[ކ�w_e��F���3�ߢA��"��%�m�(.��V���I�vf��i��bOK��^Vĸ����ѢDi"a���D�� x�$�QKo�����9�[�'o�M�:�Q_��DxS	D�"��f�Z���鲃���MyZ�� ;��\�m�z�&:�f�Qmgr���&1��onf��t7
+f���cA�=t�/���n0z�+��k���)���Ik�xN+����"��\� ���VK]޷vȢԾ�Kg��A�,>�鞦�!�W�iZ]�n/MP\ ���w�|��G�.��f�����?�len������UW�c�� ���C�ׂ����n�a5&�.O�������M�Kx�����q�aHȢ�����ԩ�=���L��\�~�/���FB%k���R��x�*r���OE�g'���.�u�VH�O�N+�'L]O���H�JǯV\��p���QX��ؐ�f)��8Z��˝��Y��\�T��~O�}�lk�=q���IxB������auӽ��2哥��~�H,�]�YRD����V�3K��%�8�4@>�q��*�Q��@�汸�"��=��Yx��ځT������R�_�6w�%���_=�7�NBo4K[E{-��F�K�:��Si��tJx��f��ƶ��0�U�[�.m���0�2�`���?�$� O��O���jn�¿��W����^K�騮S�8��xվe�_�v�SG4?����b����փ�Ҁ��wQ��fu�%���`��T P�>�����c�\be��ك�0H��G�Ǭ>^�:�-tN�nl�)_�]Z����^�t0�h~v>�HŸ���G�~��۱�hEӸ���է�F��=���:�Rw|�й!�t!��8j��-z��Fؽ�#��:��ԟ�J��u�_������I���ފ�G3����@ms�x�IUcھ޶�Р���V��-�Ǹ�~S�R��M0�eL�R��q]����Y���5YG��W�
 ��^K/V�s\/�P]��~#�ی������l�}��VNm�V-iF�r[\�cQ�f�q�3���/,��6|!�HLd_0b6t:F��ر%Q�j�s=��+���.�O$��ܣq��U�#���!��Y�,�ԓZ��y(��W�pD0�
K�8;��`'o.�25�o⪋�<�J���ZF��7����Ԓ¦p��TD�r�X���8e\�;j$~6X��z#�>���p3�Oj-��7�����A.IOL.� �E�yC�+��{'UJ��
��@��$xJ��3I�4��WÌf�(�9n�����EK�&��N����O�a����0��P5�A���uM�H�lҫI)��g�a��|�=�	S$vA�F0��mc�;�F�3�W�o���T��r�SV[`y~�L��pb\��/iQ(_�X|F^��~��}�h�Vs(ى��P���wG̰��������r���������U
�"3fh&�%fW��‴���&�_�@��q�d�Y�6e��v�#^��avD��S`�<J	)ď��!��g���Nk�-��a��R-��>��4t�(s�lK���Qt��E�|�7��%x��
Hs'�@ �v�?��C�=�͢�y�E�B��p�> �f�?�}�V�����_�IF�3�^�4G��3܅^2�4}�o�(Ő,�Xξ�6����+
�^�a�j�����{���0��|k-U�3��[Ne
�b����Ogwhg���8̂�$-QV�@!ݭ_$({��d�]ax���' ��F9W)�7�����F�{K�G ���N(�W�,�c���2�6�^��r�6%%�7w�������f���ރ�|��R'%�����yș���`X٧���:���V�t/�jo�p>��M��q::�ɶ@6
n%�<�2"YY*|�kϾ55h�-���G%���+8� ��h�k���ݽS[,Ok�1��fG��"��0���K�Z5�	��\�r�t���l�俧��.^���
�de��1	S84P��U|�9 �C�_ J��O����:����r���0:?D(��M21�,��N����/8��5 Av�1��>:d���}	��?5�a+���=~�q��J��	�ˮ��c�7���s�w�,TEZPl-U��i:B�<�3�F����h�T)���̆�އt7X`6���>��]�9�����n@�8MJ��G�������jғ�&9��@��0zN	 Vf��^��`<��d�0��Wt�Sh����C���P�}���9��j*S�#0�����)�����4}`��QbIAQ�Q�h�	��*����R�I� �Og �F
�S=��7�(����!k;p����mɗ�M����!�앵zOi����J|�|_�S}F��g!;�i�xY�ԫ��	��	�:�_&tgL@�V��"2�kԋ3�C�!E��FS(��T<(!��8{!����	����|�Ƭe�}�xR4�&��dG�~U>���D=Z����l��7m��uI�Y(С���	�" ]t�1��*�r|�0L�A4�����/:g:�l3�-�MO�\a�z�!�?L����(�ڑ<O�^�I�d��z��A��]O� ̢�ޟN����x�!HP�8�w�R��o�2�Q��R�ma.�(�S�H�� �iqG�ԭygl_>Fb����)#_�}��`�m.+)��GHV�b�#$�ݏI��*��5Ð�����R汵a�"�i�i��R(#,�S�鶑t�u.P��CyK^�Ũ	h����2��B?I!Q�����ө���&�c߼��>��fc��Vft��{�K�	���QA̒��z��.��@Q�g̮���K����䉞,�FL�@ý9���������I 2�61ޚ��ņ�m��C>+^�5&diY�'(^4I�	�{�WG<���N����څd9N�j�5��n��<�5�ؤ��
��N�����<?%����V&�3d�۪��L���v1�т���ơ�
��l�f*|�o��f���N<Q��:�z�/j�0>\�{���|�m(�;�5���y��G={
P^(��H0} /2�0�ȶ����}b�����H�nqf0%�cl�u]��|�����f���G#q�M��T6?��wA�պ��lԌ6�(�ߔW-��@SOD�E��`������O�k���#/������M��[��2�ؽ�g�oî�P���B��L2�@ ��6�<[�5A`��(��X�z��A���gl,ĩ�B,�!~Y��J�Nnz+3s���4�(��/J@���W1��(RF8^�����W��f�����S������E�P�x�6��|����VA���}��I�]֪Z@�MYU���U�xM"f���8�)<2*���B7� pm}Y��C$_^�ȿxp���I�� ���{���>	ěG��F*W�����ܺ����3�t��*"����;��I�Ёq�恾D�A�Mos�U��e��"�L��#"�*/{�����d�Ye���퐽0�&!*鉏��,7�D��;8"�ͯ�vs���\�Jť��uؼ�Z�[���5Ͼd��q����m{!�kR��4���LQck��h�t�	�'�V�����[��΢v��]-�,���n�� z��x�>\��o��_��P&�k����أ�hg���~�ַ�\�66b �PS��*<�Y�"r�9́��Dc�̐^����ś��ha_~_�J��N�jW���8��	������*�~j�NR<<kst�S�E&Ӻ!`sә�AEV��u�R9���qN��H`��:cfA:�@�p�d�pW�a�}��蛓`~���??d ���q�[�%w��3�J�`���؅�;�az�L��j�0${d.�\ ԓ�"��#z4�A�9E�Eϗ�	6�>����he0O�6>�u���7搒� ՟#ѷ�E�zāL�n�fӐ�9�i!i�e.����J6�i�l/Qo��|��^?~�_t��\�;���(���V����{x��Jݘ߃Kx<�-�/ �hcpM�A��_���t��(�J �1��pn��/
m��w�Te��+��mW�Z�i�[�x����$ϟ4'@( �O��2�i��;�IY,�km�z�*��'��aK*X��;3�W$�[F%�H��KX���p������6@�J�KG��S���y��v�h���~4ʆt��H��ӵ�_�̵���t�3dyn3����IR�N�Y6��j_	��&Y:�,�7�s��,�tH'bw�ƛ*�¯�����gϊK��^Jf�&��2#Y��p)p-@VZ{w��O<!�,�p�K��Ca3H?�*�U:湔���]T���Qv.О�|�d6d�=����+ ޻��<�h��MN6��j]<u����PtLj��{d�0i�M�k�v������5z�������v�Ƭ<Ct�TP�����kO����n1�?���bx��s�
L�#��cs*aLg��	!M:�5�.�w���m:�U�.k7y�B{���BR����%�)2�	�_�\n���Eq�x,<�mk`3���<Yݤ�t��z�ULA�:�Ԗ����3	L���c�g��,R����Y�^��/�;�����Y��|��o�CXg��Vg�U
n��^���j��v����s�K��Z��fUe�P�N��Gx����uBe��^�͖�/��p��L"W1i"�[!���L�>� ��>�l~��{1Z;B]�O��qS���Fp����7��i��U��P�[��o�ER���!�V�I�gTd�!-ȟ�k��nLA�H�֕j��Z�SC�P�'�3��\p�9R�9�EIc{{����-ߥ%�'=�ජ��z���������{jS8&I`��8Y��2���<lD�2n��#<F���vEl�����p�4�J�7=��X���O�fءxU��>�GD�0�$���V��_��	�\7۵��ť��+����;;2���{�C�gA�*���!(h(j����E�:w���ZP>Y��s�i�8����������'�a��ȡ�G�Ey�i��"��Q�����w�y����Ѻ��~tYE�Ksf.qbNd�i�i8��c�eL@	��K��\QT���p������ր�@b�l�D$d��	w��3i�.�F�"9<��w�S���~U�AQ8��I���29�~�4ݱ����Gpd�x{>��3���P�=�#��&�?f��=�#l̗A4�S4����!b�쾧QR~�g���`7�{fry�
�~��� <h�-�ю�?��������3?���*|�{n�5�X#�w�){5�Y~H:Ih�)�2���y:n�ѝB<v�-�p��j0B4�g�$�RkS�3;�c<y�cu[��҉
n����|�ԟ��o���b��tx�̭S�����M�)����QR���-!CB�rKG8��d�����m�&��sY7�6_ڍ�y���vf��ʃi�n�8Ҝ�8K!h��_\y�HX�N�~?��`�-��AV����	�iV��m�z<�]�� �S+�7�}��bN�]���B<^v��Y�|�<��q����Q-������t)�-C�j�C��:��g\�`[L2S���j��ň����0�`���A��g�ƨ�{�@�qbY��B|_�o���{>����hz�#��͠���y�^8sx�v��2����xh�K��>M�9_<a�RNåH��������>�団���
��r��Z��>�����4�j}��i}o*
9P1v:y������W�Fl�jjL��f�2��a��o�ޓ�_�^l�ϰ�m,�2���m����n�Ϳ/�0�N1�J.���\��U��e���I5���n�7��D�I�������~���p̾��!�;��1�P��4|[�kĒ�Q4�z���=Ve\�#�`?MT~F! !k�� o1wAeb��� �%ps�]����4��11�����Zv=�\�]m�K�A������C8`cO"
Vl��YNh��~�������S�l��gF�o��ՠ#����{F�[N,�������hK3��A�G��}�N/��Y��y��EI��r�7��`Y���v��s,������x�bN$S�$!=�v�BK!�"����7��rro?�J�����K#�����i�ᓣZ>��ʅ�i%hi�;f��˩��a*����Q�;:n� �o�ћ[��A*�x,���j���
���?);��p��u~��kS@���Z�`䂒��O�%���u�m���WV����}o�V��$���;Y&��\�f����PeW�� ×���cn�F;t�7�s�f�������Ǉ�A� ^�'в�W��U��[��ߴfm�+�N)�{~�K��V縀�85�D2(�ժƽ�=ӥ��1���f��I�3�B�v�LK7T/>�<�U�Y�Pa��������wb��]�M���~1q4(�E�~Jk��[�L��n�	�����.�B��Ϭ���|��<��,�l=�tQF���>H\��c�M�t	�`�1A��}�>:U�g\������LF)c�7���a�i3��y�l��Wȉ}7��[2�rV�k`��aaE�!�0����1X8 ��Pm�o}	[��S�*�7`h��U������4����f]���@+].�ٟ�����ʻvᇣC��T�nK'��K�&�)nvdp�<Fl��	q����BI9V��!is�]�U���ۙ�S��� ��������2� ʵi�me���?w���&N�yK�cmC_�HIv&��
�+��V����Epr@�f£�C)��%�c*5�;�`�s�"�}�^Awզ�	0�2	R�� &L���)�"f���
�����+d3Fo2��������g�T�D�o-�0�0B��v5���o~)�ZT}c�04Y,�m˗�{8^غok(EIR����<�oV�1�w�S[�р��Z�gv�糭�T�%�T��E�٬6�/k ���e�C4��!���Y3Q�X�)���IeЛ�)
�#f�E V�3���y�
�c[O�x��|�4b�A[����,"�^Q�֖\:���x�;���q0���>�䑂ӷn���!�7���3HRe��&#i�ε\����[��wL�g4c���,��cc�5P��[�5��d�#�8�䉟��.֘y��M���+f)���}(Hy*�J��`��Л���_pz�)\׳�NA�Ҏ�;>P���L�[5���7�2�1���?7F%��j���yY/d�s���U���K�zS�n3���%:ŏ
�xM�&#�ʠp�0F�yv~�;�5��F��ɝ ��$2ĸ0L��F��+i2.G!�p�_C���B���ḳ�Ō���p����wN�^�۞UC��ҭ�t��T��O΃�@o����jH��jv#�'U��F�>zS�uW`?��Ѡ݀/�鯂��6I��Up.����)�r���+W�1DwO����mc� ���\]�ڜ��t�bg �WsJ��_�>kڃU.��_�B7��~�:��[Ξ�:�햤!2�Ĕ�����{@.��M�A�����h$S�H�]]7��>VHw��M��Q��{�A��J,w+�PD�M���e���"���U/-�B��8/���`��
\/hY
��ywj����8Ƥs{�q��j<�o�I1��b2y�{��y;�Pq�J��m�wV�����(%��
� �Tlt�.�$fJ��y�*�Ӷ	��}:���$�s��6k�x%»��ܯ�����}��^������z�05nZ�z(�����@$�XY?;�����OM��"de��οymua���V�(ê�`�ߡ��;�r��1'�]u���`tb�g팡C���t���W��a�w'��&�UX_�h�S���,��w6Q���O��쭚����A�8�3���/q��C��8�PȺc��n�T��C�b��FTi�V@���M�Oz����X��g�b���QG,X�	��Q�T��] ��J�d�-�7�v�?�X��$��)g��u����$r�dR`àCZpv��� nW�X��
���U����[G�N@lv͑���N@=ҡ�c��XL�m��eE7��x�r�wN�2���=
ل8b��4I��-I���+&��,�	<�V4?��	K��������Ny���@�����ac�*`8XUv\A�8t�![?���G�~�B�,(�K�'"�?��A����W��e�1HФ��^�E��h��-��gJ�=�2؈z�۴\k"&�zwu��f�S��dٲ�P!c}���ڏ��[@ٟ	!��3D-:F��Y�wtu�.Oji=�?�;.�g.�'�:�5�T8���&1D���^�ӛ�C������uS�^���3�8���Lj�Q�:���i�6�����Š�1�#�|Mf3��}w���D�/2v�r��\׀�!��'�g��Ŭ��W�J# ��o�c���+�=!Z��6��_���]��(h-��m��	�Scc$���4|�)�t�b=�{."���Wrmn������]�?J������/tA�G���J¾���O����};y��	f�:2�jEhK�g6H�SA�������)�-x��	0>��i�����ٱ��d��Le}�wa�*h�˓���Y[c�&����R���]�W��� *9y��^L/��#*�+��x��I�"n�I��>�^���[����ۮ�_V������(e����|/��GY���"�*
(����I٘ŀV
����MU�(f���6��B!�:e�F��4����	|P"I$SWM?�E�T��NM�&��.2W��i�E}��zd
�����j�5.Ny��}��W�£���W�_˔��N���Pkz�0۞�1N����L��C��D�46NQ�� �.I�
�O������Ģ::8<K�v�mu��wL3}���W�o��I^Z�	�]p�j�?�h��ڰy�ˈ{Y��C��OS6�0���g�f�̝ɒ��#��A��U'��م�KVVSĞL[^���v�����hB]��n���C�)m��' Ȩ�Nd�����&��pM�?3��q�Ҿ}������,-�lU/�X�@o0���>�j�s�����G���$A<������1�t��B��X�+	�Q�RϘ6���ɏ��׈!4pc�'�T)0�l�D��������2�8W`o[α�?��Grf�`�vg�v�찔�ft�6�e{B���D�7K&aƤ��pht������� �?lM�MB��8�n颫w�����3ـ1�r��bF]�O����<�|P�4���2�?}����`�v��H5�8񵃉�M����/Ș�B!Z���54�b�>E��T�ð�~��l~�.�T�r�m}� �;��௤HO^N�WH���~R�� B<=��-��v@��&�NCPs	�K)z�,W��*�┣k9�\6�K:��L�;)И��s0�1�H
�d�P:;�G*v�����.�ݰ��ɋ[�Ԍ¼�o��E�k�v}��Mv��(��W�{�< ��c�]��h�g��p���QN���Z�#<4����ݿ{�7�Ԍ��	"P`H���y-@�c�ʹJ�C^I�N�F���7�M�Kj����%���ٳg���
=<��Z��f~ү3M�cc��S��m),ϣ�ڋe���3ļ�h!<�������OJ5R�����L+x���`1Dr`
>�������9L����th�6!�I�@!{,{�ސ�	�ma�"=�fK}D��Đ�
�3$FH�$&�$�l�7�)���.9�˲���y�9ĭ���*�1�}"��H��s�����$�0�����Sa���헴�h4K ȍ#*�����8zb�Юn��;�1~1��)	nŦ=և�o��}&H+s2�*r�Vo����+���8���x��Y�n����d�^�PVbu�ӂ��E/;R�<E������Q� ���h��^�e�J�vzcX����+�fK�/��@Z&p�r[�?�Ă�ߞ�\�7gi��e�E��O.��_����S������):�E'|�����#�(Z(q �d��CZ��y\�;�9ϼ{���N�g\]�0�� ��d����$��]��>��M��`�kd�cf$֠�1w<@�%y��Y>ӗ?��9�x���~邡��m�i)�]�4|J��X�Jp5&)�`�?0�6��!�0� �����g1tt�d���w=�QT�TW}9�Оެ�}\n�ٵ�97����q�޿�㰅�%���$�	=��f��
�BI�-(u���-$U�ϳ'X6c�9A�w�.��xc����g_�jV��h���9O��6�<]���j�F��6�w峤��O"��bh%r}z�a�o3�m����߬}�٘6�*�'�O�b�kE�lbn;b�&���S�j� 6�w�G:�pu�Jq��4 +��h<�����4���cΓ��/���������2�+�'�q�A��;V fZ7<��f<��h������.dC@����U+���~�{�N<nک r����sӬ�c%�Z�ZI�D�S��󝶮���F7z"����j������K���[������-�x��|��S���Z��6&P�A�A{oۦS`�O��Y�ߘ5�Z�`�
��?G�nMP���V(���$�e����f��_*�O��N��_��Ye�<w��	d�Ɵi�2.OS"U-��+�i��Ti^N]�:�c�9��;�Y>��4�6�ՀpG�c.wH�g#j��rh���߽�����)o ������ӛ�,�=0� �ڭ��^-�MqKv�#j���*o@�A�^:��j��pg�#��h_Y�7��� ��E�m:Ie��q�#H�<�e�A����3���.�����t����������`�|�<���j�)hC���w��æ�"�3h��ɳ��d��R�;:0wMp�<9K�6��(�A�=MH�T�����ǹ Sت��t��^�Dd.f@�F:���/r	lPԷ'z�N��H��@���8U�&}34L$�$G�w��:7�Y]�uAJ�sd����7���5��p�,��of?b�H�bd��������'��!����s�V�.�8(�;Ċ������8Mw�BP�7rts�Vg�KKjU�KJ~j���P�8ԇ������f7�45?�"������x�0u�3@����ّ,�縗*��!C��]2s �`�Z��hoP�2��:�q�����"N
���v�tP�P��č�����Sc�M�6��Z�^�B�� ~����"�`xL�����-�b��җ^_���˕�S-"ɚ��Y����j��׾� P��	jA�I,���Űer�R43����>���r�� �L~I����������_�*nn��P �<;\n���ˍ��4�R:yy����Vi#n�T��_��ʜ��ED�S���A:��/�]�Ϣ���y� �����ĂS=��EFɵ�[9�G�����R��6´��52@`����B�5����Q�XA���Č��&����a/�����h1���j'������Š�Fԩ ��~���G.z�矹����W�H�M�r�su�I���\U�m�ЬC�s.���[�א����fԀ��K����T0.�0<�^�.�bޤwEϟ��.]��I^�Ū=�Z(̦����F�}�cn&�xhA��Q�Jш��	�6)�zIG0-�f�*��@�)�l�~�\��
ݼ��8=ǯ1y�&�<n��h��������f�u��
�Ʌ^e#���������B՚'��T�6����F���N ��>f<�{Qh���X�W�g�T"�)�96>�����<#@R�r��J�ix��5�h�,�[��{��i�"­q�[�^�̑yD�e򀃙��#�n� ?���c�E6����k�1j��|��~ɬ�^R�_��P.F�Q6�CF��Iḃ���������λo��ͭ�S�=U@���]�qD%�{�n7
R8� �4�b���Lz�V�>@�G]�_P���zڝ�� 8�����ܺ���rG������t����cx��`��s<�^׶�����v�4�������o9s/ښ�[򛯧Qh��x��'��F�Qͅ��_I�4|��גQ�q6��1�e9eI��٘ �]��~�����Ub`���Sƈ>��Q��-rm�:�p�xQT�r'��r����;�*��<�D��J��m�V��QA���*n�b�)�#�����L{]�4aI����:�z��V�sW�2�4o�X�n�l*!� &|P��^@>�K��b�0jD�3�����/���N�Y�}|�������9@��\G
��P{�AS��NSlpvz��Qu��Ͱ�N>��tӷ�m>��-/gG�'N��LC-uvv��t�>L��j?�&t��x���m��	*�@?-P��i:��y�zY�q��8fc��?�OxBh���%��D揕�/��ׯ���X���3����`���i�{ KO�ı~�Ю��C%��!�⼷�͍��h&]�V����&L�x�oR�M#I?�8gKY/V�1�W4X �П�5XJph���~�7�3��S���v���rj�A��tL9���;�]	!"/#�M�%B�� �n�<��,�E�� y$˩��IK�����aFe�q&�,j�TR��I�>)F��G�V�m*�Y��&SgP�	�ah�HiX��$;�R��,zu`��&R3e�H�ƨM�'?�S�������͕)5��$`��z�0�0e-�z��N�����l6I]���1K�������un�<���`Dڃ��Y�%w�i�0�z��׋Zj�u��H�hҸ�������酮,��U�`a\+g+�6ţ��?�g��Kl�!�hg����@.�����nd5<���}���z�J]*=����O��Ӝ�,�f���/�:�p���N�͌EΜ�WNgU�r�('�;om���j��)Q�
_Y@<���X`�}�8dJ����v239"��S.�8d�������i#�э(B쁞7�0�Xfɴ3jM�n����c�Ì^|/5_�_�*�}�"���hR�.�"��G�PPz�_�s��E����,��]�F2_F�J �m���r����R���Q*��Px��K��.s� �7�3�n�K�礣�
�°Z��b���d}3�+8��9j�<$5@'��5"��x�?��mN�e��
���;�Z�gW�}rq)N��n�"״nUb���,<c�1�HT3&�ذ������O�c�����B��[����@w_I� �d ���2��*V��2'�F���e����aU%Z�0/Y��v�Ǔ%W.�(x5,���K6���K�g��*ב>?���"i3MI��4�)�I���_.'��
���(g��G��P�~Nє��r;���6��yp� �Z�����,?a[|μw�+;)��TΈ�4�����5�咨i$ֽI���op�Y��Q��^V���Sl2ak���6d��5+���������]v�e���i�1�PR���d9'i�%��V�e�$i�D4|[��&�+G,4� �a�R�
��M?#�0���{��/���N�Bfu�����vV���C���W\f̬��Lh��QV=����1R��"�Z�X�~U�#�r��B�^�-��c�n���ZG�ai�P0�Z��C�Y@�<��#���e"p9ִ�jᢁ�ږY��N����C��-�MS�!��m��z;���s <#�C�U�X\� ��"��)�)�E?�S�rY��G[�q:�W"��'��Y�0	�|W���-p,�з�9�J�E���:�g+�d��$)��1Q��K�Щx?݈{��X��TF,�ܵʦg������\I���f��[%Q�C���auUK�G� :�3e�lMӔ�(5���)�������{H'�{W�_���o��z�BgT{��
�g����H��\�Y��xA%���Pj�!3B�*�6R}�[���"���8��R%�"/1o�;�n�o���_Y��]�Џ�R�E@v���!4O4���8E�9a��V�_�+;b���G_�4��N������!���$
��5��<���Ogb�C@/B(��IK&m��Z��9Z#�yUy��U&ߝ	n��7�݆v�l:.`�����HZ���PN2W5g�2�����t��,uG7�8eBj����b$Ξ�pwI��6����Y�]��ў���7wK�k�0]��B[9���̌���)�D��_�F�"^�G�	�Sh�o7�3~P9����@�O�N����i1�E[p�>&�B{j���f)O�K� q/O+}v��[�c�G� �1��Tu������u��^S;���ܙ����UΔ�`O��|E1�jVw�2p���q�����JK�
�h��`��|�>�o��ET�4wV2�z}�u���	��I�+�$Ĭ7v�=y�nZNg#��źAw{ը�(� ��_�}��6�?F���TO��g"��0PO�	c�qe =
��K�֐�v�|({�|(����k�����t5�0Q&�i�����~�af��q���m;u���P����'�����c*�xp���z)Oq�ϱjX�L��'ZQ�(Q�`�88\���Hl�g�eg�������A����q\�pMC��瞪{��H�(��u�ԝ_P�6ﭓ��V� �393�٫ԛ�~I�R���I��L�k.�#�-���$�������f���"�= ��<���z�E�So��y�5&F"�����pȫ�>0>�p�C�9����u�mg��"�R�N�u�J�n�bq��n�+�b�u��s5������%^<�5~+��U.�Eɿ��ė4ܖ^�<�����W�rk�]��pT�#��e��ż��� �����î��:�b¦)�K��r�G�2��te�p�X�u�
�#����!�&EWi���[�1��oϿ���3�P��L{�)7������b%��'�F�L�e�=e�쭭+]m��3�AC�%�u�:��l�O� [�(��������|�R���l��c���SD��$/���OǗW.e�1��0R�$�O��b��=5�=M,U��uHV��_M���Lq��Xӵ2C<P�FFSZ�4k�)�d}Q���H>ʁ��A��ONڇ��E�!1�$O
�nZ� F���Q΀�\�.��2uj�)�s!�[{��s���G#*��[PjIe0I0Q�;.W��?��q��}��_�O)!\��0'͙_�d����d�^ۖ���4�:���ݵ���˜g�a����kΗu��y��Hw��]7���H5��
�k��, ��(_�v��vQbm��	�@j��:��>��d4#���,0m�Cc����/>�i�D
z��{�<	����ٟ�eq���'GW:��de'
��j�Ye�����W�q�_�o���lɤ`G�Us�����% ŰY�[����99���h�_�8��2�O���H`S�0�#K�E�p���-��گ�J[pWT���jc��)�4�}��9D�`��a�!��ؘUӼ�9y��h$׹W����f�֫��λއ1���'����߳��k{��*9���ʘ4��c�� �>�6r�&�we�xgI�ꋟ{H��I�Q%��w�m����ҙ���)�o�β����K��A�TR׭�� ��Zܢ��]�jv�P�B�@z#k�#��	�|W1buuJ�b�I�5�>N>�Y�mYu�����iX'>)�BZ�C6�$��J���\�dm��Y��R�f�t���	D˙Z�%:AD��$U'Q��DdT���$��m{��ۦ\���Ax ���H�}G|�H�}X�MH*���4����e��p���t)�<4|jB��S�c��/!8�İ"�:�̳QT�6G=�L��9Ȧc?�R�1
X�Iu���>JiI}cb���IZF���C�Ȗ��D�V���A"���lӌ�d
!t�� >$�K�+S+;rkw��=]ۡ��Rf���Mg SR�"�`��[�� y	'�Hؓ���|�u�Ʒ�δ�@���E9w$O̴�)Q���t��Mfͯ�R���l�'�4X�KUs��*�mWPa�M
����8*D��S�kD�3�'�Y���g�u<LI�nH�L�9���.DU<�h��n%���ߌ}V�c��8B�ح90��������\�ĥa8�]f��$����J �H��f�<V�Ë�~=r������o޹�s������ �+#�(W�t��w�B�'��7l'��R��a�>V�?���g����7�+*ȡ[a!C%��Pru��2g�H�r�:��i��-'��T�VsIH�ʏe*�v�E
ޗQ&���:��!�x�&8MP,�y��N ����Գ3�|�~]{ܵf�l&%�x�oF/���Z?H��Ƕ↢��1@��B�����P��?�_-�5w�m粎�z���r�L' (�������Q���8^�Г�zK�;�1`� ��5�ԇD���F��^��ǃ��-}V���tVf�ܓ>÷����耊�:���OB��zZ��tL=��y� +���z<ڶ�O�[KfH����âsP���T��6&���J��貌n��M8f�9:�U�f�U���Q���/��]|i�뺨m�F&C���V�ó��w���`�m֮ĥ�U=f��h|��j.�{/��j+G�����F���?l��!m�0/$��C�b��2��d�������Ȝ�zT^����첍׵�P�yĕ';5��w��d]q���}D;-�D��qA�֍��;	�(��_����|�\��G���U+�|B��x�i��.0�?XHQ�"Ԏ�BcE%
�
O)��l?��7C��*�����!V�t��xF��{�7Y62P��l�|w�P���`<�9�s�
�H�^ȧ���� ].Iu��y�c����;T���7����v���9�a� 9��� .bc�@�=���{�N�M�$|eo�d�����g��P�^E"T��[J��|�^��>�0���+���ѓ�1_P� nѸ��E�<o� >��n[��6jY���sڰd�)���S�(���s��k�-;{pi�Όڈ�l���|b%w�P�ׇKD.� q&'r�A�c�Õ(8-i ���Wp�/0L.s�9�x=�����AW�m���S��֊?GCN��ըQi� ~5��!Jt�Am�a�!>;@��8����z�1��/�RP3��e=g��>��L:�s9.��,;k@�ȶ�'�${�?0`OI����T��Tw���#X8.��/�`>x=F�6�x�`��2�<t�!IȈ�r�E�+�ݣ����X�zuђ_�E��T�u�9mN��>�E<!�O��&�7=�>��}' ����9>Σf~#7�9t"�O����vpG��w�ܷ��&b
ھ�h�I��O��̙ŏ�褭����ssum���=�F,�$�\�TХ_���C�t�9����Ǐ�YӶ׽����'����qZ�%ą�/�E��lu܈�w���h�����h��6V�x`>{K�����T��"Y@�Q$�#��0 j�k^g��4#��tp�n�T�U�^�Q�#P���R��t06!�k�u���Uf� �Ƨ�/w{��_x@�����k�^�8N%FL�Cx>�x#t(>B��3�1(�W�l��pꉆ=���'�%��A�U��N�p�	/�STN2��fׄkH� �4x��Ƀ�Ks��LjN)\��h�|-�������_�g\5�OF�)�l��n�g?oբ��xa��������!�R�,���\��\��q�� jx�Ъ�#i����E���}���f$��# X�ЩA�j�$�&`h��\����E�麣�[8�k�g��4����u������)3��O9.�
q��"X�ju")�ե]�Sh��K�D��	eqN=��m��)zu���S��q�nuת@�k�F
ቡ���[Y�L>2�H�N�ö�q��ҥ0�҇ L X��1>S&�7�0�^/�8g�����r�>f�1��io.���Xr8ّ��(:�T�o��{<���5��2iisNO��{���]�Ж%m�a�z�+�C\]y�ͭH��nOGe$|9���@󆕍ZawT{���C���G�ch}^�x�VX�n4�K�����`-R%$��dbq�y�r!������fY-=�����(�S�lM6���F�ZX�Ҕ�RPhZV����Qk�������N�0�'�*6��%7�kјeHc�=������Z��sz?��Q&\����ԙ[���ml�|׳����}�h�l��7�"n�&҃ �T�9���I��t��=��F�X���+5���+h�v��>�y�nY~K�U$:�m����R>�K�o�]�	dG�LrEݮ�ə����#iG�dx�S�%.���U[VF�P}E��[]�ORD(}r	�����w�hI������cC���9c都��,�����I�d"��ϡ�V������Gs�y�1�i�Aß�/4���`Ǖ���j8Cv��΁O����ę��\'������Z���F'��"v�]��m�kF�!�}P"����c��O(��-G�u�[
a�H��z8�]͔V�ѿ�ӂ��T6w�*��6+�������-7cЄ5W�
�P�{��f�:���0�]:�Z6�.�j0\�p��Qz2n����r���A;���!p��=��1��G���6����)�,�	Z�=���Ei4]���*��½i|����&�T�:k}ix\��KE�tH ��z;�(�	�x*/�=��70Y},�G�y� ~r�W4���U\��I��΃dLba�> ���X���<��Ѽ'm�z�ϒ0�I�'8���=��D�J�o��8vi�G?=�jo�o]���UJ�7��O��P�;�d�]�NFe���ŀ�UC_�:�D���~��B+IF	��}4w��고�Ӷ ď�k�"I����'� ���=�f�	A��q�-��?�(~o��e+Yͬ��/V�����e��0�E��1�ЫmZ�R6?�$���K�w��&;������>ӈ���'�͙\ jf-���o���K��Sͷۻ9����p��2X]g*��s������yX�6T0�>�l�������j��jM<[�}��iA�\���2+~�1�U��5j�P� `��Yך����������s2M%����F8����t�B�}���*?���bН��,w����?\b�1z�eZ��_�6�>�H=o�d��ņ�z��ٌx�.j_R����dxy?�c�߃�Z��|ty[ǚ�yڇ ω�e�e`���.ri
x�ǘЛ��h��~��d��('�07l�|] m?���!�e?� ���c@9r�{�N��7(��p/�T��v稓g����YhF�D��a)�&�Cԭ�dڅ�+��S��Ɯ���@E�s�,�g��Εԑ13�|rȍu�8B��!�PRX;g��R\�	� �&w�B ��-��̜<Jn̚HX��P<�*BvF�yK!�r[��� fA�yF.���x��v��a���KWe)��^u�A��E���.�"F9 ��t�@���O�2�/_�Y�6��˄OX�Ym�[y��W�-�� ��]�O�O�����{�ȥ1����=�;�A��O�S<�BEO@Ɗ͗A��㒫��-��{��\�ϼ�U:�W|p��8؀d�C�� ׃@�[����|�p���:�7+)7����6*+N�Q��J�Zj�Q�BhQ\���&X�M��u���
G��qe���"������b����*��U��ͅ�vC}��klO�`5�� ��,{b�ە�O�K�|�X���*F���st��j[����шΔ<�#�b�@�G�*<��{�w]e,��Ĩ��k�ȧ��9P�h�����\Q�d���x�e���]}��k�wz��)X��ϸ����e �O�^��s/F0/��2%���Dh.c�j���`@
%�L/�4����FVݥ�+����:�E�[d��W��)3�g[;W����[�ǈڿ�dAn�XTw�=|λ���3����j���`j�RǨ�f��MSVA);�@�Nl^��ff����"�����&�L���@�?��ɋP�Q]8Ƴ1�o2Cr�hoh�"7l�D��GmJ�J�Xt=�p#q�6�r�wo�Rv��T���� �ux��둼`���
Us���:��,����:�êu�ʆ,��sB�De��˥�q����fY/s�����0�O��dk!�ĵd�\�BPJ���17%.���4R&�Bw����
<i�a����a]@��鮩���R�4<�TX,x�Q,����J��-	���-1��H�<S@+�?œ�e9��2@}�a
�q��[�M8x�`ic&P�7Yݭnk�۬z�B��C��@k���,�w�m���V6Ž���[C��Vq$�����<q��	Y�<�يR@W�/в69g�0x�_���Y�M��@Fb]ZY��-��D�1\BY�|������u�1,|��ګP f�+�o;��$����;"�X<���J������
J��Ɋ)�YxQ�$`�5�/k+�|��y�6=���D^��y�ɕ%�yAJ���2� �[�@�����ѥ��:����ق��U��Br4¶nZ���-�S|�k�W�M���*Et�u���of�?N��#F�}��qK��z6R��8Ze0��\&��u�E.�X<E7�ԗa�6�y�ž�[�Q�6��%fE|�H:[o�8(!����)3�I���+_	#�m�����ό���� y�@ȹUg��b�%Q������㻅�^�Hfo]����e�tR���C4KwҨ�c�ϖY�����:����]�@��jʅ.a���~��	l�i�@��+��%m�EF0{ {x���l߁��Q3o�� �б�o��Ar���Ϭ8��5]ŋ\���!�G�3S1���
��U�SP �n_� ��7|���:}T�:�O�(�K�=����O��K��*+RQw-���T�󋴆F�G-s[���6�Βn�*QS�\fE�[�1:��8�>��l����Ն���`2HrÔ�!l"|�Ȼe9%�c�;��ݲ�!�r����~��kp�f���春W�E��"I�;r���,%ɧ��?��PE�:l1��*��d�c�Q��ø���]02d��o9}K�"	�y�e!��[��G�yu�k�ȧZ���Y�4fX����_��)�`�Z���縦���q��7�\YG��޶5'@7����% Ό�r]P�ġ��Y��&��L�Q���12��g�o�QU�C^KD�=��?����?$��`L���]v�����e'�NNU��Vje'�4�>��X�_s��)�ve�����7T����KU��!��hT]NK����Ů��`c�]�G�� H�e� כ,��ㅧ���G;��͒p��љ�I�Ts(C�� Y����B��C��T���kL��U��{�I�����w:*�k�_�� )ԙ�+���P㾼�|��kA-��e������͠�w�IS���N[cȼ������L��({���C��^Y�!��5vH?���8�{�sEk����NR��^a��m�t����'�rek����h��Z�>�쿝��
�@����� �����A�'�������t�?��!���O��O�_Br���V����w��
<�^�1�c���f��Z�a�?j��R.�~
)�˼��bTZ㈿����n���
Ən���A�������s`$���?|<D��e`�Fx�*��{��nD����,W�W�j�@�4?��I�����7��b4��!�ΤX�Y՛�\ݡ�=γ��~o�0�:م��N?q�/z�8n�ତ��b���I�\S߂Ӻl��5\ ���!>h.L�:y4�Х�R�ݟ�Dn6�k�b[ 6\~��n�c�׷2�0|�;4D�J�lӡ���g�Rb�)�[�����o.���hR'^�1��8!^�~ߛ� ΂k��!����.��`6!�#q����k2���9f�L	%FrE.R����Jѽ��Y�=ڀW.%�ܲ\NS�<�%��ӈ�ܭ�!1��k;���+�3з���M����h�{?ԍ��]��"���S%f��=������׀�����4��_�W�z0xC�x�r�9K���zH��pJ/��u��1�It/|���K���D�Y��}(ʤ!X<�M>�v۩�BWkȺs	���9��ȏ����D*�t��'q1�#i�
r�})��s�-�ǖ�r�SG(W��d�K��j��8E��53Ƥ�/��J)@Yp�I!*��ϙ���UK�0���7�Ь<�^��Ҭnz��yim�0�m8<��l<���'��!]�W���5v�U� �&je�l���{tܕ�bA>4`W�
3U����)�m|��"8��������|��(�����E��@�T��)�ЪT}�[q�)�ݯ�y��!C�j�y��nH!�b��ŏd q��<�/�>��5_�O�*���`%	3篡�W����g���+1a0:���$f�V<���`��%�}����M8��$iM7TZ�-����ڃU[��{�.a�w�tcЩa�YO(.���l�O\����Pb+�A��Q��[�(, ��YV�Y��{�*M�G����*���9^N8m0�[:��}g&ia�l1s������̔@*�hǁ�?�t2(-��M����AE�o��8����$��#���9GǓN7�'j�D��ö,��df�o�f�k�Qx�Nq&�p��>,��=��AE��������D�Z]�!i�B��x�<`�5"ێ>��)CQ�d� һG�牳-�d�~3������
�q�`m��������-�Cy{�h���6�[Ήa�tϤ�<m�
Ė�����E��6o�;�΄d]T�Dq̲N�����Ӣ�G{Ձ��]5Go��hӏ�<h��dکς�&g�U����b�*�h�4��=�7(#�8sn��6"��Vp�W���2=��؁�@1�QulD��8x*XW0�==u���ن8�[��O�H���B$����=�_��էS��9�V�D�N�*���<���5�c��oo�E�Cy̧�|�nE�XES��&�t����3H��v�#����d���|��p�D����ڔ�ʭO�������:�������n��k�8��:w�6��℻�vK���B�7Xc-�*�[��*�=v�۪R܅i�溢�����z�"�\�&^��[�?p�z�&��c�A.�yۢ��x i�����'�oov���+��� �$
���Q�)f]^8����ێ!f��$T��#�"��D�i���<�v��c\�_*ȓ�l������BӋܰc��z��G,_3�����:��#+zc:pQ��9�"Z������D�mC����2�K	��d��J'�����r(M�s����[��$龵%+���s孆�P>�Y�8��"g�P �B��KW�OQ��D`�|�����h}W�a�iWT[� ���8�O�`�#�I2J�x��3�\��ϕ:}�+��]�^�	��ܐ�`��=SDϴ�H� m5l��%~�m������"�;�#z'|Z#�Ѹk}_y�qy�9�g����+Ƣ_r�vlwqF���4)h��o9���vH�W� �|lw6�C��^>Ǆ�hlb�]I�-h�6F4����M6T���3��#Т{�����m�qw5����Q�UU#im��y�o�AT.{�YZ����K�%δZ�A�7��r�#7TA��a�ˊ�v"�A���T��,©�r?~'V�\(� #�Q<�Q��7�f��g�n���G>��X��˭�#�h�U��C��$C��r4�HAcN���Q�ĭV��}c&���sy-�#� p��5'6?3&�"�T�MU��IH��gM�{�!�_$��y�G����U��m"��;=;%^|�Nq8$�F�����k[J�A�Q�`�N��w�<��g:4�	Iɝk����ͅ)}
�f�����S��4�jkd�{���옐K�E�.�o�v�17����v&z[�f���o	%?���XI����|�[��t�rK�ծ��Ⓝ�!N`I�l8�/k	�B~]Eb�����5���Y)7��`[�1��)X������;y �D���,�ث��6�,\0Y�a;vM�Z�������Y��G0]?�Q���j�x���3�-uv���O��+�X�z��$`]��V��%��;n�*@���aa�!t~�f�y1j{fŢˍ�>�2�SX_�A���x�Қ��\j*��L�)@��6p'��8Jg\bjeEg��Z$x%���Bvkә�$�JD'a���4`M��7��dhU�O�vN��<����-��l�dO�Y*O.��9������KZX=���s%� H�B�g��I�Z������[��q�Ђ3Ӹ.�3���ڨ(8z���P� р��0�����_�D��>��1��C%I�š�j����@	R�:�|�ԣ���]}K㣳�RV�� ��u*�xY�#����K�Wȵ�wx�cxdA͜��ؒ���)ź
\ a&<�γO:���D+<vZ��x��M��������U�e�\�Tf�� �-��p���6��%|H�~���B�W-��yS<-�	� �E�>.�;�<T�yb�����bn��J��i�#��G	`�����F'{��` �$����/?1�Ĕ6�`S���ɀ£�Nn#�\��[�@|w��m�~�c��W;)�D:�w �� �!�D*ӫ�K�jT�˞���j>0�}C|��C�J��X?y3w�Px����E(&���lq�ӿ���"W �k�5*� ��R��g�z��(H���c�s�%�q�\�	XG?U�N������8�
�~����Ӓ���ъ�*|м�#�@����8�US��|ن�;_%C���Tl�N��ב�V�n�W'3Y��ғ�:�U��mv�8)N0���U�i������}\V��.
�-*��z��> �8�?pDX -�@H'A��H����#�3"B3mK#�wC��eN�A�.���i�"�=դƥ
l���
Ȩ�c5�H�I¢� �!�/1�㛒���e�4��	�*c�g/�VĂ��y;�
�)8���~�{(���J���{��bb�'L��ۄ_�3�;�f�A[�y�.f��Q����w��&�K�į=�)(�6�"O`����A��������-�+�(��$��w@jp�(�|2���8x�
�lː�fY��3���XSq
�;�U�g�G�1�3Wq2E VI���?�x;�p5m�`�U,�h;T��S^�N<.ڀO�#У�?k�Q� -st�j���'�������[J~�]�8-%��Z�ϡ��Z�Ј�L��)!�@O����"68TM��a6)��K�&;F���Z�b��倆aM��H���7�93rV_�/}T�s���Į����.=�c\��9Z��+T�F�T9����`k�!��k�z�~3��_��g�Mv�";�޶f�v������$&���x��*U.�6�Aj^�N�W��B*�ϐ���|J"� V#�a����X$Qį�]�#����gbq���RB[��@�O�#���0ٍlE�~�����i�󰷬C��Q� ���E[�aP�����N�F6������z�ôIJ}(����T�#V������S�2@��%ء��K�~��xA�h�N�������W��f8O�j�,��d,��!��L[.�2J�d�{��r���SI��#����Aɮ !5 `_,�w��=�T��W%^7.���p*�F�;΃���[��$9��P�s����P��)�}��c�g�3ƺ0�2�>����v�Y� �wIn��[F�~º����F��@1
�#,`3����.O<*�R��ϙm����b�ؔF��\�y�7띿[غȄ�=�?��HX��7�X��u�Ԗ��rX���;�^� �t�#(��}���[ �f?স�~��E�\�������wE�B7U�{3އ�~�DRN�������B��:-s�f�tG:����'W�,��4���"�����C��#�����v�� h�ի���@�o��Yղڀ��l�6;��5C���`��)�鰚	=�x��!.M���ً��g?N��yBҼ�R�?���oDf���/������%��o����ƻ�52h(A� [������R�*��\7��?n�<F<��pW(����+���CL��9i�প���M����d�3�߇�@�.�d�έ1FߦV|�Rg��+�]����6��3�f{o�~��"�b���+�����D�a6�0���:��$YtB��ܦ�0�����m*��D�2h�k��D.m�n+�%��T���έ<�}��	+�e�|�Z_���2iO��{R0vu�$x	";/��Qz^\rs�dZ��
{��a�4笁x���j����,��-zd�!xH��$���&"c,�%/�ع��h屼��ũ��<�U~*j\5���ؖ�[K4���F�������Z��zF� #��c�g����g�X���/�W���-7�@b}VIWCjZhHR"af��#8B�W°���8Hs�2V��"r|�b��hIN�ɻ�ˊ�<l`9�8P���R�f0c���+AW�T��)�UK܊j��Ԍ�U*�C!"�h ��JgC�T�|�:v&K�.��8��?_���(�D�D��	��jk	��a�A2:魻0MV��I�E_�n�Wv�Q�F����������9[w1�Q��6���"��:˚Sl��������x���d�1s�4�|��N�<Pd�	Q�A���0�s�ؤe���%|}�Qc��\�����c���ajqZ3�U��FF������	�����~)��b���{�q���@�k-�:낈��FpR_�_��O�z�(�r;VQ�˰/d��yrִ@V�:e)DD�����ܗ�n��s�w^|��o��/��hp�����V�*����|$%Exb�D�iC�H�߉r>3�. UPo�#;���4},����%ik�g ]���-}n�H�?���k^��A��y������(O��O�o����I�I艹I� �tap�z��t�������̀E�uO�evRĝ�e��wV�O���I-</��~�	�-.��K��Qm �4y�i��1����GlMNyL�dT5�֪QS�1�R{��`Ϩ���<⚧��T�*;|���,����9��#]�_�|YJ���u��<��R�r�8���9�D-əl��r�]�.
A:Ϙ9��b�^?�a��p4���b5��t��n��%�O�QՉh�]`0��]�k���>�`�.O��d_q�skY�����ſ�,�Ѿ��r��]�םc6q��+b}T�<�Cu%w��?�୫����WRF�x��N��][�1�<{�2提%ɷ�_F�ciyW�a����b��A���c����H�>{�hC}��4����8�w^_6��Nw*�8<�t�Կ��@гd�e!�{`?sn�x����;��?ԥ�{t�{R�M�21���Y�2��CH��(5v�PQ�G�=(�K�v�᠗!�g���f��_]}����ed&I�2��m��z�]��uC�9j�@�v;u��$'6�ͺ%�p�����#[,r�j��_U���~�_������4��N4�GE�jP�X<��ЏM����_l��r�(J����ȱիt�5�H�'��e���+F�gI)1�X�3v���@�5��$R� ����E�6%�Tpς��W%�1n?�j
V�%��f���u �U��7���S�gCq�}��z?	��\��rV��� Q��"��(��9�ϑ3�+`!Ҵ<�X�L�2����=,����O���ͽ� �b<�1������L�Y�8�^<2��d������UmE����H��i'G���?���8�FB@`��#iXIڤ�Yй/�����DQ�Q
�� �}Y,���HFg�M�2;�uyr8+��mo0ŗ�q�~R`Z��c������MlX���+��X��o� ]���X����|������1���.�$�.������{�z%/u��&֭[�`^$^/��8͎q^�SEή#�U�ar�n�j�)����V{�~}f����r|�;�ʨ9��`n��p#����c�v� /ه��q�6P�,�T,�f�F�Z}����/���A!`���3���B7{��?2;j���"���Q�o��-=�L��	�%�3��.:����tD�kdˇ�J��rH��&uc�HK�%��q@�^G�d֓$��~�P(���o:j��"��	��7�KV�~~���;��b})�	�_,����r3Q@'�O?�