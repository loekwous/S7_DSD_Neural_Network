��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w���N�?ƨ:�`����א"��/K��"�Bxϫ����P��n��2�]&P�V���� yx*�X*  >�5'(�3�.g�ZH��$Gn�udG��"lG��e?�6oy(�h�i52�tc˱�:ǵt��>P3����d�w��!�uY��t%�(I��������K��օ�kex[�I���&��f肼�:9F��v�6��d�x}�n9�sF�!�hH��%HI2`��"�#Dϟ�K� ����q��%q{��)yt�NhTE`�aw־���m<�P %͏�="z�Ux)]\x��&�h�1�ԔJ]�^]2�*��� ���/~e�����:����Co���Xf(n��oHU4���[�S��s������'�C��MQfI[�8���0�_l�Y�C) ��i�@� �6��R^���%y�d��)�t|���7��:��K����Jҝ�쌇]	�U�r\|.�Ϻ���7L���x��JL[卼�nP	Q���3*��V�� ms��JU#Gb$'���Ka�q�#�X�)�����oS�ف� ��X7l� ��gR{a;e��������y�ú��o������� 3�;��h�s�<V_�ߕ�0�
O�<��HN��UtފV����.6̲V_�~g�&��Vc*��I���+� wܟ�	��+��Z)��Qǟdo����n�$����|ۦxj=c���(2�W[Sh������k��o6:���v,�铦}�"�5���GTj(�7� y�����P�L��>��S)l��ldVk YM	b�41�4v+�#��yǀh��MJ{	����I�HΫ�x�`�I��^L�Ԗh��7R�i��T�}[r(ίT��Ĭl�����x႞O!��5�&�-�oK��d�vm�└�C�G��u����@�޸ߣ�O�N(�m�:��#�Ȟ����f�_.LDai�ک�ܬ����D�������u���+(�W���[�zk�O)���@��������e�7��*(�b�a�������y�P������)S^�#R�3�Z��_	*RK��Y����_��d_�)c`.G�|Q��h��ުN�x��Zg{�I}���(�� 'y�����SX<,[�i��M��<�V�E�*���zk�
�2 $l��^�D��1�dubs�6�iBI�|���O�jdfzj����»�?���C�E�!5��g��bSUx4�M>��e]��ԍ��y�.W����*�#�̥ſ��!�~/9"��57��ь�Ǻ𐷛e��5&�ؽ�C�3�b)N.�^��1�n�~��9��R+�2�
�Y�V_�8��6_d�X!8���rg��5�Ǩ �]鄜2�����(N�#e�P�]KRQk���I�;*�ծ�9��[���iт��^������	�+�$a���d��	'��|9�S$������}G�_q�Ĺ��s�8ć��p�}^�N�k}�n�'�u�p�HռL �����~�-�,X媅�]vud����L�F�;���mC����=Iu�` ����Γ�^�{�o��k�E�o���S0!�@U����}����ZC$z��A�Se��sy<�8Q��G&�n/8D�i�i�Dj�	�݅�6�h�n��Ek�����Q�?�r'J�˨�6E&ۼ����pLfč�!�� �,�
.���j�ɶd�y�h���5�;*�>E�4R3�pkl�tM��ʇ���j��ƛ1�w��ϵ��~ OL�a�Z.��I�m�p����P����h=D�V?�ҳ>1�����>���T�Rt���t�ڗw��)�vkϸ�N�yl�J�D�=�Ө�&��A?�e�͌g|ɱ�m�1}9��8�"w��S
�Q�[�b�J	x���0Ě
ҋ/�]MxEm�9��}YY�J�Ω�Īa!&�ܔ��1!ӿ]f8���~+*y퓛T�5y�j�����O7G&>��I�T9�o88�(�n�%�+�v�\'����piSS�WY�ظ�Z�w�^�߳����6�
;r�#��b�/g������#�A����3�؃�l*�&�v2t�3o������F� �Ҥ��&B@$X�t�2B'Ễ�j��LK�#��[S�}��<�̇����Bb򲍳#�'�����<��z-4"�B���u�,G�K��CίRrʁ�@�aܤv+�����U��Y<b�D��@���������x\�ƴ��[���7ҸA\�(~��#�����Oo�O�E0���Lz���w�t����!z�*hb��zaz���Ԕ?�s�<�3�yd���f\�]}H}�}Ƶ��&���gK����������yS���="�XC���/e��w��mJ�Va�Oz�&ꢇ<��r��1�V�Ӽ~Y��Fs{��>"��`���6Ā��&*�ܲ�P.����iF0)*�o>�0D`��;�"C;5!0-o�����=���i�F��zG�w�9)�����ڃ멺��x�8K��Z�	�-�.*���Ģ_����㧩���dd|�e�|���W&�9 �w�=5:=S�ϥW�&�\=c��:<��V�CF�?^�3���2�G��(l�ŭD�W�G9-_�@4W����y�J��l1�����<S� .�)�Č�g�}�p�ϰh\��d��$�\q���jK�|�۾��-[�WU/L�G�)�B�/.��-f8^U�r�dJ4H�|g'�8�CĹ^����(��rӎ):�%�"@~����E��J�rf��H�	@��o���WG��i������zco�X�"5���/x<��)��N�0�g@������^�����{<L	O?''g�@?q&
�B�KÚ燧��=�q�l�xpெVt�YsR�����4������}���ߌ*�d�1Z�SbTF�3�|d��A�Թ�<��6�M2����q��B�m.�~�"�^��S�܃�g���]�8e!�RYL�3hgUJ+&���.��/�m�o��ǵJ�;�U��L��W���!��QZܙL�/�i]+qБVt�ъ̗�Y:z|=��U�>���'W?{���|<[O�x֓������>j.�c�O�a�i��4�1�_ё@u��7޴��*�����c��@��ݨ��ʊB�dS�3w�?��ԭN2�_��V�C��s�k�̉�	��~�ʖ��b{{:'1�i�c(�9z�Ы��,\*��a<�ɰTOe���D%>N{-�
�i���?�	���i=p�H�9�j]&�!��&�zH���˦g�
����(��FP,b�נ��$���kE�5n�#�Z��5��0�؝�>�d��^���3NO^!d��3{qmR�%)���-�&m�X�K�.Q�T!d�ĆR�^�WXH���s�
��	���忇�-�Y#���Iyp�]��Qڎ��s>1Yy��F� M���Ћ�5hmr���J`����fz+5��x.m:�*-��|����[>7��6wF|\��6*z���]�0�'���Ia��n,5QZ4�G8��rEŐ��M��q�v7�i+l�ڳ��3ʋj\�靈���j��K#��݆2��;i���m� ���ܽaPK:��U����������G;3��A�K-�]�7�K�<�ȱ�"2^5�&����X7Y����2.�Q%���G��l���r��Fl6`�q�V��9�H��(y�S�QHcC��t�z2����-s	d���^n�X���T�wו���W��{%B5n9�>�訟�K#�(���H	���"|q���c@08f��J=�i���8�	!�;�u�41��|C'�\S�@�j�_L�U��\�c����2#٩:�k]��� �Q�d&��!� e)Up�O;S�2����x%fR��ٯ��ı���}}`�&y�4}�3+gyz�)K]!�U�D��A%�H0� �ҽݑ��+��
Y*oc���@?�MT�[I�TU�l4x>��6#�@��h�@�Iq��(���P��b���.��(��g�ZM_�!��	�k*�#Y�E=z
���&~�o���&��|�1���me;�ɡ�l;J+rm����	�q���HKQk�'(���������|�ސ�"�l݋�ݣ&G��S��h[�|
L�>r8N���1��Jଭ�T9���\1�4��䝉��.�Fb��Ǌ�;5ʾ��)��?�Ǽ�L�=�lב^k���mB̿0D�g�����n'=�ʖ��#��ne
(Dy��M���g���W8sם˕�v6�@ S����LȤ+/+#C,e�M��!�=D)%�2�ph��@�8)I���(��`�<�H$	�>G�&�8���2�F�wö��h��c~R�;��-��7M�l�40�W	��e�b��QL�g����q�}h�hv�^��JSTV����c�4.�]%��)������y�b�c�p�������]Y�R4y�q��=���Ԩ��9��[
;Kou��$�0�GV��0��}CU�U[;��߮QF��k���Wu|D��_^�k
���xxI��+���Fʆ��
�-��r���1L�=�f�0̔
U\�R��qv1��&�R�?�h9���ӈ/:y_���'y��r�]bf��F`�O�I}b��?
��L����A&��[�؋��l�HV��*.�H
r�0@�����lN%������e$X�D��'I�{N�I�G�i1@�W��~��q��5�=ҷ������է��1D��"5)ʘ�*�'�Q:,9�F?�>K���e�{E�c[e�K�>�!-��b�����I��-��!
�%f�6c/lȽH{��LX��`�/Ð�˪��G��FHO��&?"c�}R�*Y�!z\NxܻS��E�?�a:��Qr��h�5�~~�t�b��8�\33V�٣��ș�ж�>ߦ����޴	"�c�� �����`�^���-�9��C�z����(�s�A����r�t^c�	-��U����)<�[�^���J�F4�|\�[��<K�l�L������QА����meF���P��@؄{�v�$��Ӫ8�[�7�o�d!"_1��("lVݹ��d ���XVk�{��ҍw�3��(y�]2o`����݌��-��X`��OVWX�U�A��Rv?*I����'ߡ��!�d�������p�!�W	ai:d�1���t��v�9OC0͘���4��&p~^�.���˖R���p桼��A����� 6Zz
D/"K�f��qO��r���C�u�?kއ��'R�\;����/��A��̀w���> �љݍ�ΜVZ`/8(D�3LkjĹ�}��}��yHm
��7��#�^��&P;p�d���4�2���o]�+��#h᷺��g�Ǝ���#���s�&"I��ɾ�A1�$���[�6"�\����&�~��^�&���>30\ʏ�����8��9��O��Z��bQW+�A'���/(J�q�*c��[X2JqM��4�9���n�ߝֻ�>�- �a��T��CjHFQ��>�\-���ů�x�d�^Yv�y���z_���� 3���oH�1p������	��xOY��U .k��������D���k/ ��Z�H��EVo����}m0^Q��h�96/�:�A�GrWO]Nl,�]8c�+.]���$������b��mc�@*��rа����Ach�\��3����+���2�q��-�F�d�:�c��[�v���^�0����Z�_��9�==ۍ�DH�{[���PG8}�X�9��t�6�t��	�	�(�B�����"� {=5�8X��!r/�k����Ӌ�'������+�f2�rq���M3f˘[)��Yi�'v
I����ȪݥWt�l�]����wEۤX�-�G��p:R� 8d�d`�K����(?���$�{&(���h�Fpn0�XQ��I6�Y���� W��N�I�B�<��I8{*��<b�����U�d�z(�P�ô�N�qR1�CE��}[KAiy���O6�",����N�w8��Ҵ��ABrϊ��0OQ~����;���'6Vh����e�\���Q����I!wR�p�KTL
���)L��s �{���a�Pp[�>֧.��W�_Mݯ���݊����܀Aw�8ɵ�Z����F\�H���3��Mt�7�+�]`gkס�o�GL�P}0�#H��s/@u�x���o����S��;�?��=�޾�ƾz�O��n�B�!O�i@&|G{��5���D�)$fz��/{4�y�����9�j���Sǭ�V:#��y�\��c��2Yt���-<��ބ�D����4m�HOpaA�%p�hѹ�y�rݥ	������6|C�Q����n{�e��4�Hv^%8�01@A�}������M��,��W=M�q���'����.t��Mz^#��������w�Q� -�&��
�ʝߊ��JUX�j6C���(���!7���+�E���6�>}͔�iՌK��`u��:m��ק������m����$m��[�K�|}��+�̸�O�ç�;-�7�b�1�-���뚵S{J=���fa�oY0:���z2��J�+6�3�0_rJ��+�Tp�*U?��Q��p��VMc��K�2�
���,�6�r��V��-x'�+��)
��n��7���ԍ`�H)1z}m>'+��"��(������D�*p���<}����L6#��H���s��%r������Eކ؊[yb��#�=3�zJ�J���%�)�����ܹo�_�t�Ң������M��=BɌ;���-@�f�0\�����ͲՕy��ķ7��)��(��'�5��L(�e��hV�y,�AO%�)�{�5��v	�#�j�9��HeUU��N���7�����D�Y�:v�J�J8x��X$(��i���7�"�TN�vt���v�K�w(S�
'@�If���i`���t��%x�F�@M^e��·��C�<7y�h'��{%�T�$�}1
��pH�γo0z^嘶����ts�,�$#U��U>����[�T���̺C��>?����UM�����a'��,t��ZE�WrC�v��b�V�k8kF-ٛ�ݲ?l9����0�y9P��`,},��Qz*�j��L�I���S�4�$�+�Sحy
q�����w�|����4���2s����5_|����g�D�g��?�h����j(ޟ=����� N��%��b�ͱI��o'�i���Q�F9M�e��	��"�$��Hb���q��L*[Q�'&^��2�9��4[�,��i�~�C)��yI���Ψ��_2?���V���ߵ_g��ߤ-��a^0D�M��S�NkYs� +�}��u�Ꟗy|QcTy{�K�G
�Ц���>{��n�e�7����xw��ŕ1��*z6��i�w�r/���q�}⃾�-�����������,���������k�9����}Wc�`��tf�7��c*7f�����^��Ӹݼ�7�Gv�S%�2���vsD�k���m9	���8r	�/b�S�:f��@)4��9fyQ��$���]ygP(�ɝ5�9}����K���)~�hD����g0�?9�����x��[��d���1��8���,�SM�;��k,ƲJ��r>:4 ���4�2r�RR�O�Q尘zH;;%̐a��;[�QmL�����s3��%�v��v�`�#��z���`�r����������B�����Ơ�Iǫ���J�� ��$��6��p`�d
�<�`��Z\�� _D�r5�ϩ+%x���N���������5tw^�*�h9x络�=n����f���y2��Ǆ8������KX��������]R�4�cc!�W���D�&����p����˔�/���"L�"
y��b$�(�E�?w���4��v���}^Խۼt�L�H��nY�oe�
��R�R$��',��}�K�b�iŋJW┊��|TX�Q�1Ę�XդtT~�(�&S���c�_�T]y-S1�ݤ�J�
�T�Nv��/T�?OF�hF��=,ɐ=3��݅>V]I���1��O�n��g{�*�W��䷬]C��%��F��fb���(~��LN��M�L	�Fxb���62����q�+o4M�R�<��b�!kq�_��Q�*Xj�MU۫�!���rNta3xƻ��Y��'��h,_�/���� Ӱ�.<w�y�!#�9ђ�'�)��nb= 	�V6��ƙ���T�~Iic������K�5�t�uU�F��@G3���'%��m�%/Jm,�{={X#�ep�_�	�R���_�S����
k�Bg��IkF�juW�s�@0�����lW��^�8�cF�Qa7^�T/�THJkz�&q��Ӽ)3L� �*n�-.�,��\_��Ŋr��nE�����~u	0^5w+5]�%�&/M&�9'�jT�'�AA���:��K<kտ�)�2����z���H�a���:���0� h�?=y
�'8�C���>!?�Z��<�>�*��S�@f�V!��\�.[��x+ݸg��;b�˅��]�x�rr�o�2��K�s\h�����Hnk�۴D ;"�tCc
%���^���J8c�+��Db�.G�B�\D@��	��<|-m��f�FNw��a��o����D߆������r�\�v�ϭl7]E@K!Z�"&�9�&�1O�}���;rʀAUݍx$`�鴛C���`UkgY\#�{uL�!��|�ƻQ%�3b�H�����}!"�k���F������K#	�� ڬ�2�� w^g �1w���4�S��G5{Q6%L+z��/  ��;q�|3٤*���u�U�p�ؐ��@#!�%��d*�o'�2�i4O�S��V�?H���}�g.v��� կ�H^�yM�ꅬ������y��AR��טj�d&���m?v�+i���b�bB\2��{b�m_4փ�عN��׶]-_�A)/�j�O�~/�u�	�+�Jk՞怺���H���8��Q�E�����y��MKFW�QiYQ�P����}�@�L{�:4�i�Sk�q������1	F���'z�w;� �b�����gVZ#�$မ;o����ll?} '�jQ�C8�ڑ')!����}�hn~"���\}�l��m��&��l�(:b�,1��i�wu�L��R�`�?�Y᜵#�F$���9�J|0��\�( ��9e"�JZ�N2��%��'��Z�N˯��8�*��X[�S���{�F�cHG����e'������P����E�ja���^	�賵�e�m�y,�����Jh��G��Hh���P��2H��>�ߨ���넇���Me4���pޅ�6I3
}c�RQ��W�X�t�����Ia� �mg�W�]i��w�s�d��!��)�0'���)8�����ty`�Hy迆ƅZƜ%Z��Ю�z��د&��l�/�˄4���9�p�����h��\I��G���(�%��3��B��9F��jY3n�fj���u$�3�=tgxD�Eڲ�_�)do��ĔY�Zj�QX����b�����H?�B� �/����'`$�%1t���Bō6�R�Qrl��k�
�.��=�p�ʸ���O�$ڧƝ�~F����p,��IoS���]�⤥���3�0��bKW��r�@�ĭ>YG�|@�o̦�s�֙��{��\D�Ч|�����X�㔄,�g��].V�;��Ays�U�|S_�o�}C��`#;X�u���6�[��& �_֒{�aCq2����>+��,�{�M����Z�D<�Wk��t�;z��c�t���>y9����[q��l�Y_G\��4/�Db͗�9-�S{(��E��S>&F�j����=��l3����U��#���h���O�'v�[)��l�<�q,]X	� :���/�_y����G$�:��W�c��)F@���uSRu���,�ѕ8}�d���GL<u|B��uU\�8Kv1Vz^:v�C����dN���6[|]��È)�F��Č�d�@i볠������3f$����&�C(
k�̣6���!��D��p������z>fn���F�u�)s����9��Е����$�{%qr�QM?8�q���O67��AxJ��q��=��v]�vdvW�e����[js3-��4d?���Ʈ/�N�'xS��BF0?��"=���m�h�;/�CJTA='	�E3,��h��\�܆u�$�$����3nO ��p��'����h�F�\��g�ֱ�_����Sk�8��\� z/�Ӌ;EdDj�󼇀cl��Z���/���o��g�Uې��tc{a��#�R��4B����
ԞV"���6�m�),�
Ȍ�Nb��-_�V�����9�K�1�R+ߏg�6^�&\`(��7ɱ���?� ���k8�̈�%|B�+������:�T1����R֛REOoJ�f��r�g6���<
�3��%�zt"����L��ȡ��/�p�����N��|U�)!;���y�fm�b��q��)j���Gd�+���*Dkʔ@��Ara	�x�m�B�d�WJ7�l���7����?��J.�P�@��1�D$M~M�*i�О����>��ѭ;:�a5�p�&�G���<S �8�-���	�������TM�A�F��f=o0D"j�a���̗�K�]�{�V�Yi|!�j���>$`1����p���[�|.��L�<Pzxք���*���/K����������{B^�����==�Ӎ��:0q�V?�������W��Es�
�l��?�Iz�� FNE\���c�+���̵���I�Q[=F�i�D+K�yϷ�ӏ��7��8�5�kr��I�