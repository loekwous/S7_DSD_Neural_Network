��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w�6V�%{�(��ԣ���*J�@�������c8Z�D�b?�;�߼�_��Y�	8�(���7 {��T&�D$o�6�{ �|D����9�R�:���?r�&P��Cf�ͨ/�ou7����Hҍ=HK�3Q+�{�#T�t�
*����j5G�9�9C$)�����a��^�Cݱ�F�實��Ɠ����׹9@e'*3Iک��ܦ�:�Z�Xᑣ0�oGC>mmd��A�!���9�*ߞaS�j��$�rUO(���Oc��w
b�ۡdX@���4nMH�3���T�),v�n>�~�)�%�H�U�M[��NN���{$_�PN`���.bR��{�#�ʃ��J�Zٞ���;��k2��F�~�M��\v����̱�w7��O��[��j�	7?8u6 �v"�FaO7�r����0���Z_9����%�t�HF�}�>�����;d�t��=����a�
�Y&jV":�����j��:���ܩJ=���U��~�-�)�@��7+��jG9����(;�A�����#6�Wo�I��P��%�r�����:`a!F�cNI�&͈e��7hq�T�Д*��7�a�=�U?-�6>�4���me!LՇ�����kh�\�<���j�������iM%��tNX�T	s -��J>��;�ʌT�\����O�x
�A(��.��d���S �*#����V�(k? ���c�*c;�B�0���ч=N�2bx����A�����i����4��ʵ�J�5k8&�k�j�G�p��A]�ߖ�d�dg2�1z<� ����?��,v4��^v�X������oD������n����g�I r�.��>������Z��W��`��QIn׫F}���~�Q�x���c�t�3750~�&g���R;x���粯#���A�4o? ��3j�T�3�ئ+b"	�����#��m�������dZ����D���::�*T��Ns �[�T�lo����r�V�b��viB�n����7%���F-�0w/��Rt��&�!~P��?I�'{b~q϶dt9΍���H|��]1օ��GS�jM���qW��m��RI�@N����1��#��&$�rj�x��* [؈G���t|�+h �#VΘX�Ɔ]�)�s[���w��6�%��m(��Q�����W��G»Hl���I��b�XB�������9��x�]�zT�6^.)T�@tF	��<��{Q�)���,h��1<KJO,�d�ߖ�r�im��H3"�)�g�I��C���²I���ǈ����BNo$�צ�vaeְ�h�s�����&p4T�?u���� ;�2�tf��˷LK��RԻ@�Y�zK��wu!Y^-؃U>�������6��g�A�'�X�#���A�U>�z�Yk0Op�;�Ha�N�tQ�5�mO��#2/PwЦ��к�_�s����J*o3\�Y�%Ekg�mx:�m��^U�� UL3t��A�� 7J�$TSPQ
�trZ���D#+�*k�I8!X�uD�u�
G;�r-��%x��Kh	���ǝIF�?Ï�l�k�ݸ87
6����<o�=8��S����!R]�,XI�sV�<��x�5���n��פ��`�"�P�o�3�I��ù��h{>�۬}J�`���¨nvݪk�M��&�tXݏ��HL�D��ʛ�8�
�Sj�/Dw�������d�\�42,E� �
14⤏nSk��;)�ι��%Ƒ7jTeH(�����4����} 78V�������?LV9���|�����6'.$�ג�5[���/g��� �9
,ԋ������a c�qBf���ֆ���R�GP#5�bנ9K��Y�|m�B�Z)��|Q6?jg��[��t5
fWp�E"�}Y���5r��*z-?��:ɇ6c�q)�S�ĵL80 �7�]�~~���R)�@�Q���ؘֈ��ܫm��\�Y���P.N����/ja��к����n4�K �X����*ǜ�/��������&��Fx_��ɓ���hkZ�T�jM��1J*��+nC�ؒ�=ђ1����|F����5��v~W5Ug��TB,Pض+��D�a�),�ݛ]I=	<m�V׾�k'��I�\K��=:u���<jES�W�b$�I%��R9����.'tK>߾�P���V�� r���t5�6�����l���J!<AaTA�}=���!����nN7_|(2y�r6�+�B�'�:�Ty(���?� �]�r�Z�+m����B�]�x�8{+2��h�1��N�)Q��[%Q������B�ɽ���DH7+�fwl�S���$�c��	�9�P����=���$���8���#��\�{�\��E��� ����lq�GcV�<�0��r���Z����/gaM����ᶽ<�!�����O�vew
7|<t*�H\9�K�TKO�z���W
8�<�[���J�ɟ��y�s�3i(����H�<aE�-_#pV�D�s�=��g���k��O��/c$e�c�Uͦ��,�m��b�9�&���<�9��`@fD__���%��v_yz� ��=�B"��� S#���m�fy8Rǿ����J�-�����h�}�HJ(���m��A��C����:Д}�!Ǐ;�[�Ȫ=���h3+��4E�kk�8W.�h��~;�aj2? ��߻�w=Fc[����yc�%웉Qk`��H	��E!ʚ2^�s
	ű<@ �s�LWPm�>T��I�F�cb+��P5�����.$�{7�J�A��Wm�P���!���l	w
i�?�\�M�JDҧ(�^sg���WG;���O�^�?�a�T������I��0?�+���6����W�\��9�D��B�n����9�Ѝ��x���ԗ ���p�چ���ڪ)�a��Y�娞9cj�P3��GD���g6	FͽaAk�`��L��vK��Q5��0�S����S�=~�����n�Uum@3@K�>��g�<��X(��yۃ�L��l����#m!���� �)GV�I����"ַdL[��u���e V� �Q��!����P�hw�)"���q|�ҫ��$�ϋ�C���^��Soe�#r%�b'[l�=Ԣ��+At^��#��&Qn�9��g�.�Ӷ����3���.�	���r���D�������R�Oҳ���IK�:W|�vw���$��|��9On���\E]��mM���\.���-�b��>ˇEE@���&K�����{YGt5SRX֌pl���P��QB����Ӵ���T>&�i�mD�:�9G\*��;���{�޲1��G��w\�٘��V�}�\��Y4`��� ��PNJ ��DC%NL8����_�R#P0He��z��O�fY�����E�^×Jyk��ݔm;x� 4+[��V�~�H�z_E�w
�*��R�?���0T�s۸Ǹy1;��N��
V�fGu�qʓ�gdj�Y8Yx�E[37BX|�>A*؆��n)��� ��E���7Մ����g �4�Yt �k�%:m���=�lqwǭ����>F�9X�z�0_@�ݡ^AW���������e�Q�!Z���v��$�:���7π�jXN��|]G|���	wԮ�j�q�$����C��
.#�?\U9���wp)l7,�Z�AΊ͏��e�=�8=�F�M�g���騖��N�;�����m�1��-���'-&�V�?F&%��b��5%������#>��>Z��U���ձ�oø7��K��j�[�?���I��5R��$���Rʬ�T�R�u�%��\m�U��~�����+�<S�VH�b����K��<s�$��&�1��hB�*io�w�i:�#U/�%���,)�\!5A-�/���<8[p��核�1%���a��EN�F[s����g�"���i��&B���t~֖W���DF5u�:Y �w�i�/�D�pge8U�=@.z������OR��W���i��P�\[B�`?�-t���=��<��\�}��GGf�`;��O���B���X��Ԅj���kx��yW���"�(�������@��
S��?8뱲�s�B5���ާ���"���	4Go�D`��({�W����1�8W;9q�� ��Al>���%ԥ�YzƯݔ��{���"��Wip���~��Y;�e.+�I�������%w��RG+�ς��A��MB8rs���>��%d�ls:��) ;�ҙ�������ْx#U��t�U�<Ɠ�_�Sp^�z(E�ǽ�F�rgK �p��z��Ėhb���z�a����7BM����n��U��G�(;߹�p��N�f��"���>I�{�L�(�����2�u9D`�����OD֓�R��A�+=�@!��Ȟ�d���{g`��.��7j����?ձV�n�G���I��~���_�Ɋ�f��Ⳝ�z�ȕ	x�U�7�?�D��S�ŗ�&���_��=��R���y�/�B�V�#�AL(3��'* �'�d�}�����~/B��`ձ�J���vt.�g��Vv��K��@�dW�)�|���a�+b��c���x]��f��-�.s��V���WA��]�U���g�Hw��z殅 �#^�52�� MQ�<_|^��l��	3/�m�����Z��W�N�!H}2�Z�ǐ�Z��J"ָ�,��B8�ك�M�q�r���j���KG� �ߚ���3��(��!*S�9�-��am�d7<ź��G�Ѩ�}��₀
���w����~�`���^��g^䢰��<djo�o�d� �$�C���&�2�u�P���":��p�
�X)����h(�{hC��t���.XuȮ��#��D�I��LE�?r۸���[���:q�����C[����j.W��U!�P���-��0
�������5Q'�lP�����*�Tw���v�p5��x��Y'Ӈ���nU�}�f���~�j��
��C%��,��j�q����=��W+]�!�e$6����H�0���r/�<�����qZnm�g+�wGX.�+�r�O����jBg܁�N�U�R9�c�����c��,6Ǯ_�i�B+%�g��%����έ�p�����ݽ�H���Hku#^Z�u��|a����z�\�(A�λB��LD����W�*DR��^�oݯ��5�� �"�H!7�_dI��(:��VFL��q�bq?���l��Lw�7H4���6�R���fL1`K��1$T�� �Y1�	1p=%hj����5����e���JN��Vʨ+���*G�ay�0*�O�i��:�,��<|�U�s
W,��N��SQw�qlT@����w[�WEL�g%� �Z��ڵ��'GI�/�q����WdeA�E>�
�\�P0�We�w��!K�^�<y�Ҁvz�Ѕ�:b[8�)���;��Ĕ��b��ʓPk��/b��ؗb�-V��Y�sp��`����%�%�D��%����T��s�ج��=�g��6.�>6	G�Q�Ue$�(�$�(jn��w&_
DN�t������t��]�-h֣��=���s0��$�3�H��O� 2���u�`6o�lI%���j���}�C��Y-�H����{h�ɼ������M:h��y�3�5v	o�Ï���E(�A$�u����,����|	;E�>�W�]�k�-���]����{�^��A��`{?%(�(�K���"���"��RO����c�";��k*����{��e<��kJ�2����H�ǈ��^��uY��>+��Ľr�xU��]���o�R�2��2F��\���$�Y�C��Z܇N�p
��=Ap���N�<09�'sR6��*�Î+�wK���d�g�~������ \z�	/+Kf����;��rʐ4(7#j��{��F�b� �g��_v��� f;��؊,y��ǖaMu\'��>�c��g߫����~f�>�x�GBt���=<�@���b�-0%(۫�TR�_���T���ʷH�cIƚ9�}�oN8Ӓx�Z��^	��*6��A�KMM28���>�M��ޅ,D���u�F��ġ��x��=�����]wm��/t	��%oЦ�rF-��l�2��Uwoڌ��g��?�� ������8�����y#c��~��$%JQ��`��| �5��~a�4{d�oht��W�ĢaNd��7WV7���ƽ<=�"x�OѺ��dX�k���C�J��YJ�9���&����E�|��q)s���å>ݷ�u�� :R\%�_�B�795p��u�U�x�[Ґ��.�����G�Bc�5��7|1vr�I\���|f������oZ�X`)߃� m�4��g�Q��8��e��ۘK�:���ʅ���3���������SzJG9�)H*oњ	��B�N�V��9ш��$��$C{7h��Mn>�.�R�GJ�{�?q.�� ���͋�u�Ъ_A�cT<{��@K�$����3;�ߤ�G��Ș��
!L�J�4�B�A?5{B]RP(���n�<Bގ�t�E�kY�/ٗ��<lyv�غ��B?����ކ����m�o	+ʘ�l� �[T���j[gZt�<��hǵ#� �Ǻ^N)N&�k��:&���,���AІ�a�M���zZw_Wk�&��n1
��p���?����沐\tXwҰ(�Y��&��# ����>�as�P�a&)%�@�U�C3̓�&0���;��b�I�ʊ��dP�
ڒ�Rp4�1�x�^�@�/����9$��]�{WRE(�⤺�v��TJQ���'�[<��F���t!�ɯO�`;,ʰ�T� ����0��p�4�ƥ�N?@!tv��U�&n��%@t�C����̦pi�o�k76�i5⏂ӬB29��̔+J�ޟw���W����j��z�u��_�������C->;j��'&޴�+qX`ؼ2	����¶�%�3�{ۿ~�����֧MF���������kr+r�?�M�3��K���^��D2���V#5�m{��Ėz��ٙ��+��n/�𝋭q������>]�6��G~m�{d�=��G4ջ{�$ՠ����"�}��/�i��e@�_�/��[�v#��~���c���K�Nu�ڵ��`A�����E�+tˢ*�Y���G�'R��s�k�[�8 }���{Mr�U�?e��i����gw��1h���>74����B�̡��V'f��d2��ű$���wr�l�P"f@x�4�w��<⺓�N�M��چ������ﺟ�=�@mfiM�ڨbY�)�`����c;`k��]�{�)X��ɂѢOf1���<��ք�,f���(<��uOg����8�_�P�u���&0�3
���p����c*��1?`&n=�����G�撞������c.u��~�BG�M��ԯP��"m���,G�zQXQ6��8�Jn�3Wj	��ݿ<��=HR.�0}��W���R>(�(���8�h�kAfQ�*���36ۂ�.F[�}�۩�{'��/�|�����ڷ����XoLU�_5Q �<����{���˫������R�
���J�����ft��d����6�J/�ݲ�|m��zf~/��(��t��N�Ɖ$����w-���:�%��b��.i�{5޿[y,G�o����Hr���x�L3f�Y�ӄWWأ��頯��"��(]���p� @��gm�� DvJu���Ɖa�(�ĕY��R�{����09�D�l��%9�6��oM�]�v���\>���|�o�q����+�*�ko�|ӌ�@[�$��:Ք�N��!��5�6�������k�~���*WٚX�0E�#�;Ztj�D]�����~i��c��ov%�đN�qƱ��|�ͤJf��=�����ȝ!�J���K(V*��4 �9�
.L�y'H������z8����;ڟ�E&=@��V�rC�m|Iy.9�1Y��N�������Y���l� �ҢZ��a44d,�j
c��2��3�'���V�f����~�yM�UJ�0""Jp��8���z�6�����ֺl�Q��w�*��#�b9�'�2u�x}Bj����������t=�4��3�ò��%��%ֶ��U�x������4�_b�r�ٚ��q�z���o�4%-���=8�>���?��!�3���ő�8@�r�-7�襵���#`����
|���d�0I�+�Z�Pe.�L�bu�rh�<t�	�X�&HB\���WӴ�ezWB���Ǌ�����AF?�����Ӕ�Ж�6&�f���fx�Ǉ��:||C�梽U���K�2����s+���OȑWg���@6k�m�,x���ʄf�a�(��a�l�7�A4|u�B��K���}2=EI�X��	U�D'�'=�{��?�u�S蹲�c{qC���g3��
��Bc`so�#/8(�k긱q%{?�PPUM�0\�����q���֕?�VYa墙5!9�s�peMJX�r�Kd(nWB0�3�+���e\�Oc<�,�2�?�Gh�c���ç.�����L�iY,�u_��NɅ�zE~h�?�<	7UW
�;�Z��.�w�E���\E����#�/Fyf��AHr����BAD���d^߹��,�B�0hN+���K�_�ɰ�'�:C(�
�$%J�q>s��YZ\2Y��o`K�z����0��>k��W�/���z*49?���G]s.��rW})S�[�{������l�]=G���r��ޑ�O����]�.�3�}.�yn�	���)��jO���cş������)-g�;S`7w���g&���ݓ�S�[�'��"F�;�i�][B��m2���\�������옩_,����m���V����Ot�	�b��8�w�I�<��x",��=EA�M��]�ҶDB��宙j�O��/1��]���Ni�Gu'���_���I��؟��U�v��VrR^ެ���A�T��T��VX����+�R/��/��-��w�;H��#j"�-�����}�)��E��]���Wr�Y~3'��v����6������7q�J�Ca���[���3�g|Ь���FF6�*R��/����ҁ��Ε�\��;�=��Ģ���G:�'�7
R/�2H��~<�8�|����2c��F�h8*A;�:b���q��"�{r1��uN�^���׫i.]=��qJ���np���a�,��;��|㨦e�38<�;q�fX�����Uw�H@H���l��>亇�֪���8��bY.KY����I,m��#���4�U��׶���C�����UΘģ-����H��i�v�Yz��+�N�.\�o������ՒȁJ�9������g�t%;��&��I�eAbVk�205,%> ����e���1��|�g��k�b��1���ahl�7Z����K����_Nk��M�{��4�О�C�d�Ĥ�G�fS�:�G�<�Kj������.����D�^��I��&Q�	q]�C��J�����+��.=��c�L�Ps#-j�� ��<��gX-�Z֝��H�tw�@7�be(����_4��lNSe���?
M���J�<�+G	)���(Ԅ�|��'��w�EO�&��B;7��5����RSl�`���l�`�{��_��Д��B�>	/����Wf�f4�|�X2^����W�[�c��2	"�o��q�:0"��Gt�q�Q+)sֹ�˭���ߪ./��|�ﳻ�����q=���^��]z�7�nm�ߥU��ë��/o΅U>�?\�7���Q8j�3U#���v���!�Ѹz��
��+�a$U����bh��Y:��j��mw���g,1�����A�'��wy�^���<6Y��f�( �[m̉Ň������j��-	aؿ|g[��8s&������&8�t6�LA�RD�~cx�㮂���������NUKB���D�0�T��@��#��ZJ����n[��������rr�T��X۔%�I��5�Smn�}�p�6����8�w7*�/�>֭f*�����'|�KD�ǟ d�-1�{۩^� �������H����n���$�����<����� �@}��g]|r��]ʋv��~;��pf���x�Y)����9��p8�mƫ��B��?�#߂q�'��k�Nb��8W�	���<
���w��)�ff	@�w�crU���hu$,�Y��7�Õ��&��������Y��{� ���B�K������j~�{GF^K�ϱ�����FL)z���;k��Bc�ґ������9�V4ӇJ�23�)����[n����壌�,��:^s����b�"7�ɟ�j���[��%�S�Ӫ��H_���$6��~G+����hY�6�s�"�	�ۧ4�h�������6=�k0>���RaИC8��GLAx[���G�'Wn	�#eQ�OZ͋�K�B�ԑD����H���M5�~c�J1b@}Κ�I����$H�WjQ���ǫ@<�������(a����}:�QS�}*�����BkX���F^��>fO��H�ye1]�����]��.��1m�=Ԣ�|A��ڑ+ʲv��	Z�˷�RpJX�l�8ċ��P�'6�
M�غ��i�8�V�� Qc��z��k������k�ɔ�E$�X���T�G>.]��LK�cx`,a&]H�`�+��GﰇO:A��X�h9��E@�%TYu�Ŋ�H'����V�����ӯ항<,��%5�w]�BE)�� l���*׳���Y�Db��=j43A���;�^>%aZ�pz��X2�L;׹YvG�X�a��Y�պ �:����Θ/[�1Ge�V�.����I--�0o�U�*�u�;�*�+u���Lҧ	��H�0�</�)�1�o+b�[w�u6*��ĵ%����;nwzKrZr+�l?��$�A�g�L��9u�&+Mt��FԜ3�.��5'ӧ�<��{�\�r�~��yd�j���`���eyО�VR���Q��� �� ��j�X����:݁
#��:n�]�^���Low�oza:\@[d�q��k�Z�Խ6�<
�^�i��F��#��hdYґ~A�F���XVۿ����bʐ��W�dU�."O�v&��TXF�Z����{��&�s]�(�.�3����ԗ�L5�ت�QI���B���f�ܾu����\�O��8��6ۄD?���6e�)�ñ�3~�f�,�I�K��Ԥg��.��Zk��o�^����'�Ga�k�����g~m��eT>3��E���z�����~auo0F��ǆg��Gb��d�ab�/���|�ۮW���Xm'�h[Y�N�w����]�Tq	 {�lVp�ɯw��L��A��	!�\��+��@�YE~��B��|�=G�m�tΒF���O�4��]����� ZX��P&��s0�� ��V�����V��ܚ�wA�GP��?���ʡ=�I��B9;�a;В�����?sMƢ:�h�H1���W����-厛�"d�7I n���a�v���*ի�`�噉�4r�|�[h����՚���H��(�����M�A�Bi��1c�K��y��q��¶s�͒�E�J�'����ꔲeB�^c,0�2ʷ-��}�)f	3}_�_��S�����_�u�8����D�x�=��Ƕw�}�f�� ��f��^���ϸ�uZ�D!|4������o���kZ�~��m��v�ڥ��1�a�����,��"Yr�f�iyeCԌ  �i����iW�5����4(4�+6�E$�?@!<����W	j���Q���n�R.SiFrt�@���d�QE��"d����y�(.�~:/��E���Y���`�(��%<�k��c��ɡ͙!���� ]��qHt7a�D���&^����p�_��[���aR���o���R[�d�T�˦�9V���f���1r�������3q���1��������ah������8�(�U0���!{�"g_������9�)s'Hu��lA���Z����Qő���:Cf˃�B���,<[8��܊M��F젧��Ab{�8�P#�$,���`2I���,�s�n>�g �}�ꑻ>zL�fW*�?RyK��z��Tn��5'��A*���7Xٗ�0���qh�$��%� J�2x9�/������(�z���?e�˖!�|P����sͿ��c�@?W�VJ�G���7�M9*?l]��\l�/�L>[<�|�a��{��~QJ��K>e��׫r�v�왫�3Bv�yop�e�'M��Vî�iOb�jѿYa��=ο}�]A�(����9��橗�{��pR�h�x�W� #���?�Y���wp�d\s$�FW�D��8u�w<oi.l{&���%�+o̸�+�7³Xꞟ��0���7��V>�ޣ&q�a��&�`n��|���{�����g)' d�Y�ՖNw�*a@�9rY��2�41/��J�`��婻��y��>+�؃0�Q5��4P�2Ba�w���` �\����)x{.��G��r^��'�S�`��S��j��E���7hM��*�V�RS�s(<S$z-�����dL_%�l���>y���d�%x�}�_l��Z���t� �r]��S�t���D·0��rmrL���8X��
�\��+:Z�@�S�X�9<X�	S!-E���j�ޘ��$��k��Z�Ĵ���7M����8�t�A��G���R��aъKd=J+C��:g��ܵQT
� m4�p� ���8g]�� �,2:8"� di�p��ޱ��w��� �y{'���L����flq�;��E`�~�Y���Q+B�惍�!G}wũS��[�pa?H
��̞3 �&���e)n��<���W�`�Z�[��3
�:7��������^�Uyz����يŢC�͌�㠑������m�J{�=H\؝]�y��P�O����Q��2\r w�C3�U�Ĩ̯f� z��{��W��y��kD�L��b�S�br��&�(���ҟ��*Έ���=$`᦮���
����:���q�2�(B���J0%��!�8 �]18$��ر3�Pr������z���h�f�s��m_3].�}հ��"D�ψfB��b�@��;$-�tY~��_�º�o�քkw�a�5�����c�-ꮚ�{�-K��\ԉ�ё:I��`+��ط�N���l�#X�#�'.���ᘤW���D�Y�5���,[�ʫ9���ϱ(���6�Sݺ��d�i� 3�k���`zÜՕ�{�.�_#{&W�Iǹ��E�_�ԑB�r� �*�(ױ�1O��Q��wn�����N���=�b�6'���5�5���_>����u�H�����@�Q9��T���x�G)��+�d&���r��~�sN�0a�m�lTf���Z���u�?��-O���3	����<��K��T�3 ��'�&���D�[��]�����6m�v�~B�l^�cD�P�-�_�ARY�@����Q�7JDc��?��EUI�S-��)�FZ8�9��9txt\H������� �������m�3����Ҙ;Y����L[qR�⤄~j�!8����qC����7�wԍ��4c�W�i-�\�O��<��& g��k��\f"�NW�$-���g��4����k)+�@��UL�?��97�vV��kW*��7�T?���ՃP��*�S5os�Nx�R����xMI��xU,�T^{�h�Y@��@�H'T����;�J��� ����}C:�0n3d\n)��R���J0a���>+|�i;<wC��U��b�f�P����� �zɟ�Z���/R�̎��5�UO{e�X�-l[���b��ȇQ�^&r=s�m�����v�Q�V��E81JkF��m�Jo�_�)���0ƫ��x�dH��^�.�$֔́���_o|�%�&�*߁2��-���6�vb/p���T��a�:�eɒ����dUi��۔�Rlt�VJC`��e��I��/�i#�'��M�^A�Q�fZ����r���^{��5�sp�	�j&-�$ԝ��;�fj������>�
ZXl��d���	��Ϊcޫ�5�j�(L���jT�f����rX����D;�cz�Rϴ�����5��[4 pҎ�N�$0�aqt�L+�I��\��P�\y�=�VJ�����b��g���N���b��Z)SD"oԖک��� ���УD��M�!F ���%(���s����n.#wo��誙 �}�=%���cR��b�&W_�����x���Ud�D�뿍��QVe@"��>/_��6���&���<��}A'�1����1CF.@�)����)y�.�()/>\��x�:+�b����w걾�n�N�1�3@ΧB��_?ҏ�&O����D\
��T�U2-��Q�M��x��(�����X#G���!��e��م�m���L3���&�	Kr�g�xD���H��9������R�fu���<X-2�;�2��E��R��ni�2��P�F����8LA�b2zP>?O._r龜Ȑnj�	�]0\��*���+%R��T��oK�\'�3��o���紉X
�Չ��E�8V辝�ԮZ���m���CS�#8|�:o���B��\�̸�(�}����v1���Z<�g����"���n<��g�+��m|Z�#u��x�e��b4�W%%�7iMʠ���{>KP�+Q���YM@�}�;�g�	�=��8���h(?V�wuv��bMs:��kd~���(5es.���z0�0h����~�g��C�����_�R�]w�$6(���lzN_'E���T��o ��w�`N���]9n^*����;=�1�áp:zC����u7\$LT�n����Z4|�&��
��.`�0�P�E���m	4��ވ�4��ˊ����ec��>�F-�f����q���{g�+Ԅ�ּ��mf�X޿DF�k�~15OX����#c�7}�4�t��
�3S�p%�bm�ܪ8��$S�U�n�z�AKB����H'�Y�]0����z���
Y���]a���9���I�^F��	��|?�c��Ck�q����[z�_Q�&LF��R=������$M�o!�g)\�7X�(�; �vS�K,�%>;x]�6#��'x����F'N�#�&��]���|����d�*�rM���E�T�٩�yw��	��2�#��ח�����3��'�ڦ���ٻ�n�8Y3�����_�oA��R�z�����kR����[Z§��/(hW�i~�fk��jo쨊�G�l�ӑ?-}�v|� g�Ã� �E����Y�xQ�H��^�����Jf����N���i�B�>{�\N��}��U��A�"�OҜRp�~�m��-�a���^��OX^�/uV.��|�����Ea�����Άptl�:��Je���EJhR��Α^,����-^}q�:���/Ļ9�jc=d�9��eiu2Ƽ����:$)=����;YQ��LF�l���B�Q�ܫQ��L��)�Y�F�Ѹ�.q����[m𭬲ó��V�X�+J�Om���#9KGT�-GP[DQ�e22���sw� 9n5AC�� �/Z�
��`O�| a-��=���U5����*?~�&���,`���~����ִ��W:_z`M@b�?��\�Z�@ӹm}������jk�_����˪Y��?ۍ�a�#�Q��n`�6�yt���'n9³�rD4���sfjuF�F��5��ɋ9M,���"GE*Ϙި:S�UR���vLJV�%&��n�)�� ���������2.�(8s@�E��Jms筗�{��M�9ۺ V'�g���?��+/�4�ZT!!�il����X��K�'�w2�,�,�g�:%�Ifc��P	̚����tf ���8��}�f�nC b����t��4W<W��6NS���0��N�6�6��i�%T��sT���B	��P/x6ɯ����_w��4Z�;Ş
��7�(�G8�����U�����Fz�Zk;
�z˺*:��m5)�n�I�"N���1���`[*�l�ղOںW{���@`[��貛ʴ��t�!Uܲ�9_$�Q$�t��>�`͊R;g�����d:#���U��z:pa#+��7BM��QJ��]N!�gc�
�a�k�~���9��U�>��mܗY�-�YŽvM���cmD������-N�9	�X5�� YhJ�6�u'뫱�ȁ�����(u	UZG�����-ڴ+8�Z�zxp1��!D��)2��;u�_5j����E@x��) ���?��/o2bXYl�h�^��x���%�g߃TNFU�XW����c-�񹽴��'��?��W�����e�.��>��A�e�.�<���b�����"���	�w��PQT�R6��jM�4�񟕦�*n�M�	F�]����4�H����а�`4�����Z� w�v����J�չ�R��A�T�~�9���wɔR��H[��H�0! T<#5W��~@���p[�}��(�Q&�[J!�/w{�z�Ş���,��OL��)�x��=viw� c �m�� �UR.��f��+��#?KHO��[Xt�����Qm��%��ݰ!~���S� ��o�_M�k���)�rr� Oc�"�u�k��P����B$���%���<l: ��@�h�P���2�V,�:��gh�2��H7x���s���L0���e��b��*������d�bF�<�f̈́�O�}�~ ��H���o�(�@C��2�WP���'�g�8Nvm�a��q��\��s$�N#&�����Π�n�deC="��ŁC�ԋ�~�7�S�D�kO�,�$��q7ӸF3�������.���K�^�%���J�^�O���:�Q��$^���Tj��p�/cSk�����;O�D3�fj�|��o��Ң(��ml�	�>9�R=k@ ҆k5?�*���u43���y���t�_����o��)Lrs�����~��V���Q÷2B~)9QIk�2�w�����1E��2Հmà6�G)b (�m�M��d��g���;�1k�~6��^��JO����9����ἵ3�#S���w�LgՐ�ύB<C���\�-��C�yD�KhM�:��� 6���{MёX�����\]��q�36s6Ъ�D<0-��
B^�lw�8�"��+Dc����@�rlm�+�3H%�B�Ұ<!͗��Ƿ���jX�j�����m��8�Dܐ�T2�3,z�˩�c�~�%¼a�ڃs�`�,�l�1J:�YN������7c���,�8���~D�b�>�s�b[<$T���96�1�����/�a(wi�>�ku����6��\���[É�xI���C�0��Np����vf��3[
�PR�Yt�*����/V,��!;XC��kC;B<�g���¯/v�#Q].f�T�*2�����,=�C$0@��UG�%�#�]����9����ˈ׷H�]���V
�B!c�o��i�.��3�,B�B�ȶ���rj���f]�/e�ۣ�Z�vlY��GL������<ΐ�s���,�K��ݸJ���*Qq�\#0�Wk�����p�vTf����r��"/vL������$3'�a2z�v�o�l؋O3�e�lfi��|��ֿ��d���������dY+�Ȯ��!,Rd��U�<p�@��!�d=`�%L>�m����D'G���y�.��f�����v���ٙ%dMd�!>��zɇ}Z�v�� $ 7���W�;��FX� ��oPĴ�]���u�տ#"̽j.��VY�nj=ol�i����#W}��Y'u�pl����"I���F��l\W�_�4S�ɂ�� ]��[���k歀k��g\a:&�3	ir~�P�֜�%�I�?�+sUJ���h&��{Go[������M����jw���xT��D0;�G#(z-�{L+�?� ����E f^��ҟ;궖��y{v�>hb�d ��raNyg���w5�5E�g��q[�R߅��d�(�$-�t�vWv�Ö��Vp�!|�DkL��E���Ƈq$e��g-�eF�mޟE,���^��vl:E����!��X*+G7ML�����e��� _l>B�ܞ�B�l�6�����,��e?�s"\Uu^����Q�t�H�i*#f�)���{�$�̏�k��˹k�~�X䘻���Tb@�����x��ٿe�$�?ں0�a�^�bm�S&R�� &$1£��
?c[q�'Pڎw�q�����6p�C���}S�u:O��7�X��&ϋ�/�z;��U�a�X=��n�h������iJ��{��k]nb�*E�G���=:_ ��N@�#����f�;Ps��I�QJd��4&���c1.?�l�����C`.�L����N�$0����G(�@�¹~ěPJ��QǄ��f Lv�9i��^J$�t_�i��PsN�&������<� Ä�X�����!f��7(�� 6A��X�,Ml�)����AzqF����-�j��N����o�����AD�}h�!&A`GT#{���*6"��7�^� �i��2s��&����eI=&(�}+�	�[Iy�>嚯0���(���~����v�5�`��e͆y����q9�t`�+2�ŋ��q��W�A[:%#@���vߣ��V�e���`�=�]������<0t���|���H�&:r�S.��AF��G��pL�ݻ��jPr�ը��\YB��������E���U"1���/�����!�¡TV�ξ�Ϭm��E����y��)�ӗ�E���PL'���b�}6FY�/���V�%P�U��$ �y%�j�bn�mw�Q}��+���؅�1�զ���귨朂,�����:���5�^٭�������E�/|1�jtd3���-��������|�Ǵ�P,��gC Ʒz;�|����cM(Lx����w����}6>O�r8NyL��PP3^IU�[%#����Ơ5�A���c�h���e������D��Wæ�W�uU�t�4T3�+���Ǎn(j������`A������
���W�If�>�Uk园������#2�h�������U�\�n-��T[#�� 	��"(�d��Nۭ�!,�9c.��w���#�?*�%�Q��_��GWA�,K˛�Ͻ�
	�gҿp��cS#�2������������ˆ�?릑�����W�3V�!X�(�,��:��p<�eB���α��p���g����2Zs�N����F�%Ѡ��Br�)U��7����;��Ӄ%�01P3���&���
"��c�b�|	��������~56��q�x[�ԞU�o7$��������!�t�l�r�.�w��/w�s�fz��I\��!�ѧe� >�{V�C���=!���z��p�ĜyV���f!���J�WX�, ��׮���a,�Ojz����o����ԃ$�-z���*�\�)���3�wH9�u)x�����)J*f��NXk���h, �/(�V���'z�+���}�Wbh�%I�̾I�2�h���:�^�B�I\��g�ܵ
����s�K�+�fY��G���i���:�M�Ɓ����vD�BQUH�d|��u��Q�,���m;Vᕾxi�Of#�e��� �Y5$��>he����%ɍ��e�1��+�ȳq7���:ouD�d;� 	�KGaE�H�p&:��2�y�D2|��Fd�iQ[��΃jȑ���a�F��R2��?G��~
��l���v�OC����Ŀrב��#�� ���V�ru}'��8<G��7ᒽq���8͹�����Y�MM+<2��MΙ���1�{��9�Ӳ	��	� �p�Vn⡔p�W(?�90�T��4^ӓ�U�RP0$��j����޷�u�5���pg&,~��s���{���%�b8�S,/h�G��˾.y��D�?�r�:!~~<��+>�p��A�������=���Z�I.D���wGNj��L_�n1^��ز�"t�O�g��b���#�C�b��RW�����RAHE
�% Ë��r��^A��ω��//|zl>L���_�Y'��s�R[�ⶠ�o�J�!z��~^��Re_�~<�m�Q�l	MsZC�D[]�	v�L��h��l9�J�_@Q	H�Xx���U�h���R�I|���=SB�����£Ųi��p�L d�&|-��H �'��5�.Y��n_��g��{����F�B����Xͣ�
9����'��(ca9�0�w���P� X�ʯI��	R�Y�F[��,K���n���g�=a�щ���
ŌO��j�ǒa�$&�(H�h\�'O�W����$h}�{<RؽQ�V�)@�AJ1�̱Fx`v��Υ�����2�uVr ��hb!�(���i�u^���-�a���hSd�[;]���݊4C*|�s�KU&� K�֏ "�A׍��F � �jh�@A������!��vsC�6����p�^r�~ҹ���Yg�}��60@Q�����D^Ƶ>�$T ���}֊�Y*�"���ڨI$�|�
��ޒ��~���拾P�Kᲃ��H:@۾����6ǽ0F�^M���dY�Tq
G�x�?�x+��M��_2
Z�*]���4\�Q��|�;���q�E���l���lv Hݲ#Z\g=�q9N9�-*�9Ԕ=�C��r���������q���)v4�@��	�N����K3��n��}�!od�!� �4�̅M��18��\���o�Jl�G�V�VCu���R+1�9�_'�	���  �Jˮ ��c~{a�A�(�����|��佭C��ώ�]b� 2E;���u�_L��+O�6�:y@Mw��%����s�0b�i�x��t�v�j� �*4�x9TC������J%[S-�|$2��V����)~Dw�"$��i���1�JW���H?I~� �ov����$b��>���*81��p�7a�ne�Ɲ��T�RV�J˴�����DG��ʁ��u�ʡ��bE����hh47�į�<�FW�6��� ��1a+�k&����6�q:(�C�8����'����n�Aƅ�NύMI����br�a˱�K�v[ج���u9U��Yi$�<r!��ՄXt�(+�%��8צ���6���H��xCu��-����Î�}�$IM�f�:8�]h��;
y�T��ශ3�~,r�m�ՁJݣT:ty����n��'$�f�9~�h:�ڣl����^a����i:e1b�NE|Z�_��!'��cX�H����)~؄њ�8����b�����Y;y���?Bb8Q�G4�������J�
�hV"q��W�n@��0B�ghW���y�?���bQ��;�����x+_[�-�=���JQ��`��"yH��c�6�e��)ȣ-<��r��iK�=�kJ
���O"�;a��Ѿ�^��7`0�<��cWk��`G�,���� ɋ0�i�N��A)��4��	)�r��� ��85��I������g5U`�մ��$���pv,78�LNh����\��!I�U�����1��+7�u�a�^rS�;�wQ��������b	��&��2n��Ӆ�����e��|�IvoCE�Q=���aZˌ`?.`rn{�:>�}�~u^G{w���e�c��+��Є.�`����J�
�9+���䘿��}K���`�В 5[�@�mk<N�VC�9�e��n�m��o��������u���>Uv
��a
i����Sy�h��XA=jc�5A;r �xM������l�S����5�!�Qg>�y�g�̡���Ҥyz��V��Y"�����\��0a� �Hܰ#��W�cʉ�|L���
�n��ɾ\p��ʦ,XH����4��Z5�=Tv����� 2�B��3�-�����
X��?��%��=g��RɾkL;��s�0�b
���B3h=��F�ϓ۪̈́����ۙm�_��Y��eR�����sg{���f��J�S�u*އ5$t�4�x���D�>�pR(��D"wQ���@}F�E��fvg��Lq0�"���˯K=��W�V5�X�!:�}郍�8������0s�qZUah$��7^��Q�M�a�~�Rt����M�acHW��Ա�E;I�aA|��ַ����}�}���<�=��sPC/=7��:�GL���u�߁�l�L��KD3����,|���$�=�Ԓ��7�\)8]���O�&�s�k����'�U� 	4{�i�����x���8���|���
X�|)�;�v7
r�Ƈ��Qʱ�R�(=�ޘ�/__���9�1i�&�4���������r�>F��X$]�*:��8v����������si3+
p�.��=oT�� �_�3��H%���qp:Xi@6�����H��l����XD�n u�����^�<<���;��S����@I"�n+��zg�[&r9e��������Ctk����^�fؽ��jf���C�B�_� �^FfX��*O���:�3����2��Z+zE0�o�c���:�`��k���Н��F�+�����%�Q>�2;ڟ������#��-�{���a?����/�֪*F������ϧ��$����q,���\=���f°y�X�?�eA���q
U;�mr��)��vUY����#��h�ء�Q&GZ����Ma�-�Άia?���e4�ꗕ|ft´��Tل#E6�X�&�S3�+�B���/�D"��Bm<"ƥ|��'�@�ۮt�L0�c+ɫiژz� B�}�,��^��L޽i:�)Q�mr8�8]�2��f�D���.�ЉC�	e�ٻ�8����T�H�������dRau@��Q	��-8�
ͼ�����g�טɨ����r�,�W�y�i{�x8;�
�J)����|�ˉ),�f��f\]u깈�<`��O(�ԷJ�<s4���}]�}��8���
#!��|_Jc�,�v_{ۍ#q����0�����WyT�d���Z�t���JB~ӂ s��^�`��.�ԟ�ڻ�$!y�A�{ri�� �������Ԣ��&��a�e�8��0Yit"ґ{��F#8:�0L����ߠ�/���є��d�lp~�T�,���u�ߏ3�L8����LI�����6z�(���L��3�i���&�D�y�a5��X�o=�ؑ8�L*�H�w8�Lq�\�X�KA�瀞��e����Z������GZva��Bf�kK`G�iCQ����r�-)�Y���M��gږ�gm(VD�~gԹ��Ό.?K�??�P��w�B�B�_���FIث! ̏��`���"�P͓�gU2|�k���\}�w�A���8L�>�k'PwkEd��T#����n���ʚO-ʡ_p��Ԝ�`�%���4T#�������)��� �a3�-�C�}�y/��cL�a��)���n=�,�Ơ͜�igͤb���tHd�J�^�4(�;�8 ��6�P&XN��.
�)2���u�-�8�����py�fS0�#0�clK��u�s<v��q��Wg6��b��#>}:*ǃ�5�j������k�˾c�Z���v�6�	� ��0!=e�?�� ,������btā8�>T�����󜆊I�8�@);�yc��`(��M��|�>�>A)���f�<%&�	 h��2�s�Aghe�}�dg��5p{WZ�Q,�@�MY��hz0�BS�2���fq|zW]����ͱ���|h�t��_�7j3�3:À�g�"���g�L�`D�̏�����`�������f�I�:�Bi�`Umb��[[ �������*�$/>��6��{�n�w�E��Fm�~�ʽ0Z�0���>Ci�8��O�����i��3��4���51��,#�@��u�EZ���l��a��9� �)t�7���>��>��a�-�t�З+~�j������=:p�2�s��]p�CB*�;�!0?�����GQ���%�+X�Rʐ��t�����&�!7�u�2���V+�H.6����;շnL���2~��.C�Z�X�GNt+� �&���cI�.�`G�ie�)Ԭk���#����\hJl�|J�9o�@	��KgԌ1�1 TO�Ub��^�J���.ז���t����*z	9�	���=��&��d�p��m�����}��ڞ{n[�0��g2%�� 2ݏ5�6�˒��Uv䇻��z#�� �A�e"޷�Z���TQ�A"Q�D5���֬F��S�Ģ�yHs��QJ3�t+V�7��2r�3H^��t[����[�f�b8�)���zt;�vm	gj�	b��kH���h��%X��]��KP����l���,bL�N�����n�@g烣���d�C���n�xɄ�s����Ec1/�"CP��p̲�l��	
=""-!p7�Sn"e۲��c� ��69/�`C�g>�i�$�h@JGn��դ2Ι�L0V~7<����&Y+�v��mTls��{k�p�1���^h�~�&�������!���7��	X�"hu$ߍc�I��X�߯[��L���{k������sa�β�+���<?gC�a$���%���RJ� K|	E��e�������6Vr�����G���v2�~}�]?Ru��i�<9����p�	Z�%̓�!��K;$��7s�����G�/P� �f��e
��AI.�����&�o+-�cSE�-��|�����(;�)�cݳƏ1�٦�?��c�\;F=Fփ8��oT;#�ʵ� �-��v��E̡*�-ĉgq���'��q�#��}g�E�/0��C�ӽ����Q�a%������zr��)�%#�;���I��o�JT�t�~�)wa�^��m�G}�3����fU܇�ݽ�j§I���X}����ZJ�����e]���L񥁢G�oT��y����3� �yv������us|J����+�[J��܍�uϸiشj���?i���O��9�xd����
-uCt(�炣����eX��S��S�v���)��)&um>w��=�G��,�	bآI~�4&
�J�*�
����k���j����T����Q?��A46��� Nv��$�` ����=h�.��r��"�%�縢�p����>��*���D�R���s㥟���q�nD��r1�
��<\��f����]<tv0$���r��5�	��^?ǶQ���ErjV�Bߛ�� d*=�s�}p�����TW\=�7k}`ܔ�t��3u&�7�#����C�M�9f�9ZV�W7��]1��\[���V{��̨E&P��}��aܤo�{���ft|0�����N�C�=�7lŝ>���o�ǌϸ<M/�,N��k��zy9�9��B;QS�rvs�U71��Z�Al/����7+f��� �3�fa/�m]�ި��m#��"���/��j��[M(�7��
O�4 ��~�9���v��#3(�%�ʽ�h�O�{�9_W$=�ʞ����S��^�:w�)NY�#*j�̥#@�Ɇ���`�z�Qо�Lvm���d�{A�a�2\�+���(
VC�]y^X��|��I_�[e?��k5��):�z.ЭZ9�7��||pκv�[�qI
ݍ7��oQW�V�d���[�rISQQ�c�������J(���+�x>�z����M�$n{"��m��2�'��w�8��M��j���}���	vό�>X��%�5xE`�����"��M}u�*<੄�ٱ�S�/�;}�?ܕ�a�is�����r!���uGl����vˡ��
{���ө����P�y���_:�c3D+p/�`!�˝_�$
�M'�H-�@��z�CAXt!;w�����X_�rB0����zq�@�r��	�- ��)�W-�zyJ��U:Ϫ/��.9q��뎋�"���Y��̾Eo��t��R�T�vnH����p�/T��0�v�}�����m�E+=�S)���bW���#��5�i��͆���C�6!�uʌJ�3����$U��u�����R��8.7F��Ǿ�z,�֮�~�����!M1H|�}\%0�Ĩ�t���I[�Ob��Eh��@&/ۖ����
T��ޒ��ƢTKV��n�z�5 �ɋ����+��"N����9��5V}�8�b�yհF9mLL?��4̗�[��`+Eҿ�mIogA O%<�u�4���Q�F�����>=�
̭�$��h�h�={_јI_�W��G'�,R鈻��e��..*��{���D�i�d16�"��ٸ"��)L��bZ3��#�3�g�-��Y�Je�c�լA}�?��� �űa���<����*^�?��ﰖ,cH���p���L�&��6�����͑�[�u�L!�b�uJ��M����VD���x!����6��l&�rJ�u�3Y�rl������'���̿h֔n�����k���>� TT�M�����Oiڐ�	�L:z�}���@��}Ze�q�6�ֆ�V~�o����p�{�[K����=k�Kf���-�2�rZ�����{���ȠOC��ʚ��?���ug���ΘZ���4>�