��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�l�(���q�a��8`K�nz�w�V��� P�����"��l��p��2����}�iH��i�k��4'�����C�H-�%����c����ݮ�ƒ/L�o ��RD\���m#Ө���������tw��NA5b�7���ßS����2�+�X~듮K> �1p��M���%���|�8)�"���*q����E�x�-k��A��#����a 0�Ԗ~0Ghg�`,�i|v`����b���I���g �2|���KϦ�}U�+��t�qYBy"R�>D���tx܂�O3(�C�*U%f�[i��V�o���W�R�ѽ�	��Ǹ�L�8hG�]Ii��o�hk=t��zkC\V�P�0�{{M�^<	E�	��!G�I��E��/2T
�qd��HלgҚ������W�o/?Ґ���J|9�4��(:�zX	f���M_���j�)F���|�M+M+�D�j�eB=GF#�`FSF7�M��լ.|v��Ub��r[>?x��IOʕb�����5��X )�^k���q�����'̄�ThC|����Z�F)PjO�X�$4�G$sH~�u�c�p�������}y\V���Ծ!s�ċ��e7�p3)�c���H�V�,�+s����v��1$R�g���x��3	����tD���3E�[wI�P�t���5���#�8*`x�����=�m��e�)�B�gB�S\6��m��'<��#���bta2��[�9n gilZsk���8�S:SE��$P'j�������wM�X��]B�o[����xM%��T�$���f�_#�������~ϛdEچG����rR�_L�˯oƓX���n�&9n�I!���R�F<x��k{=*�fٹX�<K##pp��]�)~���'��Jt��_��zR�l��M4��9%x{���j�X��A;w~Z��^(qp�:�wL���?�L����$_����rWnK��.�?
�nc�M�w�ȍ]�о��·��\���M�+����j����ԋ���Pr
�����V�����?M����W�v�ȩv}��T�Aq��lx�L��� �q�O��ϐK7٠�_��만9���[�ç���^�.H��E\�W�p�� ��C.i=����-5F���c�+>�~K7��=�}�ڧ���_^������7� OҾ6DIX�%9��X;���]���bec���6Յ|!��d<��J���]X(N�U��A&��G�z�?�R�o>�F[�[5)T5ߕ��Z ]�:�����8���5A���v�<�y�#���o�^t�8fbA�ٷYT�74eP8��ZUe�/9��׎k43��ӓO�b��0<М-��ua�(3D;������.Cy��XlT�]�+9 ��&k��j��q+�^�Ϛ8{cd`5�<�Ǉ��<@��pu�!�.��z��|,���o$�zʍ�c:
JN5�O��6�{�ڇV���=�ֈ��0,���<�s���E���ȵ=�~��	U�B�ܲ����_Z�A\���LS,����� _˸��f�누�z��-��Ϸ����(� �zi�r`��t��$=�^t����S۷���º\ N���
~6X	���^Q�j�Q���e ��?ӾIMN����u�n112|�=7���̫��&��� Ax�F#����HZ��x����B�\}�t�Ocs�֮֒A'��n�ZG�[�my�t �V�&���\>�J릨�"�he���ߝ3s���)L��坪��4�o���s�"����[�Da,hB��wA�0EK�*pF.Q�J��{���Y�2����V���T��R)6��y�=5��|�^C�$P��s)/Z~�]r��2�-���:��ө�b��'`sr�/u�M�MK#�dF�o���4���{��#�x��e��w��7��*������bW��msu��OV(yn��QG��(�FS���`��֍�7B!�fo����޿�t�0cǷS��a�9H�-���#��|�9>=S��h
+�YnN��E]1Ʒ}"�1�><&ٞ$�SZ~��K�L{�$�譅�<LJ��>!V�碟��t#��� �\���G��e2Z`��3R/��E,Ɯ���{����F����`���,@�M�nw�-�	��P�	����.�������b�\)y��e���=�.Z���3j�^}	gϏ���4���F����$\��D�pL��󰯭���2" vz}�ĿA}&���(��_5�n;z�����t��m�F���f/��ez���N�2_c�Ӭ���1G����o�$��+묇mz߭�,(�7Cyb8 �j]����b V�r/�ǂ��=��������{��a@}>�@O��-^�[9~��X�}%���u��Ų`g�!�q����1���(�[�ë����2�:=�ᥧFh���\v��G\��k�f�qr�������v��S�i�E�����e�p�׮�]�}әL��4W��<�kO��V���WX2ryU��x�jʅc��U'��CƩ�L
O{��Qqf���?w�@=F�޼=���0��_�ЯO��n3��d��J3����q�#=�2}�h�M��z�q=e\l�־U�J1	�f\?0o)���6B!ɢP��/˹�t��.��̭��M����V�g���J]�C�1� ze'��[<��Mֺ���	H���o$B�X2��-����m����zҞ�G���`�%YF�̓�H�Ζ>ľ%W��8�U���Ɗ=�"�4�ּ��ۦ^���������3W��v>�G��#��ɿ�"M`��[uyЈ���Rȋ����i �0�ETq�RE~<mU�U(N�m7`�gT�Z�{�m��T�+��i![�mh9O���aB�%�Avp�x�Y�?M�t=�{i����t�BH�ߑ^�k#�H�<TKP�%9��p=ߨ[|hM�Yc��g[�����)[��-��'m���j?�CḺc倚�ɒ%�v1�����#ڸ�v6t4�'�?���nL���<��nn��߶"��lk�����Tx��dL��3r�u����H�gf�l;��w1cB�QGc���킫��z���o��K�D�[ީ�uɖK��c��|��4����E{E�D�@�����s�\s���+q��w/+���Θ����7��?k�VI߮�GX��2�!�03��ù}z4���#��2K:�B�!���_�R�qp-d�ϟ���C���w�n�����0�~��� ��#X8��f=�T�z#^�w��A�o�6!�	CV�B��f��4(Kc�1�{T�w�Y:��=��&������%�M�� �μ�W�GMn��ד�&���Li�:=�H~|W�M�����Ρ-i<�z���g�gh�����@r �N�T;k�(K��P�/���穹���̂�YΪȅ��a9��4�;��bzɵ������V�DL?~�Z��77�����O���V���U�w���d��+����s��M�<�u[��	�ـ3��w��  ���<���e}�y_�2����%l�Q�m�"B�ǰquus�l!�)�5�����]e��r-�����U~�V���L�5:��
�8�3�
��H���y<+ :�u]&���K$��l%o
�KVt]����x���6�Mp�'{�Ck�$BB6�$!�:���w7��U��,�)��K5��J�*j���x�E��^��#Y�-WY_�KN�h�/�t0^ -`��"+U	Ğ�Ɯc�ӛ�K�N�f�b��|G�������R�M^�&��W����:N���g�~���'��N��e�٠k�#.���uA�'��S���͓M���k��Mr.I��Gw�������,��G���m��*�Y��T��E{�Z�Z���H��1�d�}��5;�tNlH0�X7"�-�{���|7n��_H>Iŧ���p�J��6խP*[�Yf��c5�Eyy���(2�:��#r�~��;'�5�VIq�LSJQK���N��A�DGă�e��i���/�x��#���A��nV�5���j��^Pڭ d���k
�^�9:����^�q>���@$ϯ�W��g%�w�_4�����&o���ዦ���J��٤�:cL�*)�D(�YVN��?�H�$�v�jq_q0�z����r��f	��7l��S!02� �D	���KKcY-�im��O�p�y���\i�48B3��%(��������_�E�h�2T�љ��ˍ��b�N���(�����o^��3�$`8�}
�o#����O5�:0�H����t�@�'�8����H'�ҪxXܞ�fN��<��W������A�צ)���u�oYqGF����Y��z�J=�$�u�v}���v^�i�ǆ٨��N ����Ip9�]�J2��cjb��ށ��GM����]B=�Es��_�M&����	C�`�k� ƾ	sp�yҤ�܌ KD �'��}}�W^�<>�I�C�׎g�gK���l�"Qz�h.b�cL�n��Uc��o![�Z՞�7��<���W����e�8���'�:L������m��]���L0�-C%M\�%�	�{I���7>Y����$~�"�=. JK��Ѐ����8�Hp	4�a������b��#�f�$spAL�GQ�Y~�nɛ*�����8�%��XӺ_�n-�#�����F�pD��L��2�H�z�&|��_����c@�I�:��W�;#z�$Jl���Z�D*����T�'�$_�/�U)���vV�q]n�$X�~ ]�(h�y�"l�b�z���z���,Ї�OB�C�s�4%CnUP_+K�t���\�2�}��%���p-%�����D�Vq̜k'lؿ�����1�UA`�-�I}-��aӬ/���r�:�vjaL��U�Q�#�p�p�%l�2���i�XBH��$E�6�#l��!`����;���$<B����!M��a߀mŰ~fB�Ks�F���~��;�Ns�4��q;�'z��|���N����* \�<�+rf�ZЏ��*�Hד�=qu)�� ?�ǻ��ǲGE�J#�;Um8�򹠔e��Ht~(nb��'d&�U��7�mP'�	���/wv�y9Un8����
��s��NC�H�����uG�v/�%t@~��	7�1�-D�Ό�M�@dޜq6��w	��*����ssѭU��ոz�I� {���F7Z��'A�D�Ւ����U9��+�Į��c%���z~ ����+jօ�?��]�X���Z]l@�C`���y�����t�-lή�+����簝ަn[���l�v�@i:��z*���W�z�Y�(toz�^t��v���.�Մ^NbQ��3���]m�==�`b���5a��;�Y�s�O�B��b1Yst��j)ϲZe_\�f�`����"�ڵQ,�Wrd=�p���s�F8s��-�_���\1�9��DK_~�2�l� +cEo�Vv�f�8��Jv���Ĵ���i!�Wc�������:�>�P��nX^��G�4u�ʼhY"l�Q�[}jm.���O��d������.��E6O{���"��g�Ċ��˶2b�;qTYջ��;TR������;���ZIvD0jB�l˨L����kN��y��#��m��87�'ޤ�[�%���~��/l�GY��O�xSg�4�ygYI����g훠~����
���[��虚��;6,��<�e��jW��a�G1Z ��q�n��֞HcS��0CɌ�@�ɖ	/6�-�ƈ���]�꯭;e����x��#�Ɖu��/�FV�t�!~y�fBvJ4G�i����;��z�ރ���{T�.�W
&ZW�P����ŝ.v%H;m�{qRN�8�:?�Y a1oMS��5pu R����4�`ʩH�2>q�|�%��s�+Q.V�t��Eߔ��$�Ҍ��X
�����d��jD�}��.�t2=��I�0(�e�:�Tݸ��rT���;I.�L���y��]b�C߽[<c����
2�h*Q'���yX����\n�Pu��ɦ��g���A+��H�F{����͟�ef9�>��R�:��wO��\���Wf��{�ֈ�\���A���]�B�ٹb%P���aN����I�CZ�Ǡ�8U��9� r��A!vXi�_8}�V�z��׵d4���`������L��@��Β��jg�n��-���,��A�E�y��s���PA�Z��;x !oP���wv����t7>4W�"4hX����˯�%����>��L�'2�ޫ��
9���(&2�Ģ�3� pnI��@�p�_v�D"-ZVe�"<�y��R9�iN/&�����2d�܁*a�{��<����ie.�j,����K6<��\ �����# ���`Yy��t>�MxZ�#��˕��t���S~�l0��q�7m����~髬�nifQ4��_�d(~��}VpL$g����E��E�z�We�孢�}�����x{�B�qNx�Q�������RJ�~�RM��ܞ%��I�9�t���ǻb��C6 W����Bm�jr�O�����w�ؔ9�j5��z<�sk�2���lw��)�b}�}GK"ѹ�C�d���W�\ȫ��o��H@$<�A�{���x��x��Qc���]k�%�^��(�ؽ����h�eH�� �\B^%�f�;'`��
vEv,�[w�<����#�W��<OC�bYח~5B6=����)��(���):=���O2�R�U�����4�&l�-[\m���g��ɿ�ꉂ�?�\�t����p9nV ��C�h)�fv&�M��`q^�7t-/L��/@�%�{<��ǉb�u7m7X�x�	�k6��g-�Q�0������x+��+>�I�Q���O%!��LE�3Yl�xd܏"2���H��>Y9���?4Ǡ�����&:�����h������f�"��&i�4\U0"ƀ�?ĉ�'��k��XĪ��Р�:�Z!���va�/�߭]����� s4�K���� k�����R�3��4z
����vI��KV�eܪ���L		��3�Oq�2Wa~�ޫl*ո�#�`�/���#����z����JJ �xp��(�c�Jw �s��._{ C<:{X�]��^P�g����yvu�9�띑����r���&��O�5n!,
����.��{BF�6d��!3��)c��ySa��|���C��/��[� �&Z�v��h�f��(*0���9"��M��	�!�<�gO]]�tה�[�G8��7����b��w�|�Wr��(��AKįz�\H��UW�[��_�辘�~��~;��@5����c�m?_|G��y8��5B���).\"���d���&�,6�o�R���W�i�"���~y����v�������o���!��� �E���K��e<k�ʮW�X�l�:�S���	FW��w[lAJC����6�W��z��%W@ez�<�=�+qEpf���Z��%����8���Y�=qDd+R�~s������|���w�E!�"<����1�
�4�xHi�.���:�MVA<� fͬ����k2�^,���6�4'&��؂<��-���"ǐ3�x�&	~�Lp��{q��b�ڲ\�f*"��Z���M�H��C���0#.�C�
��bv�&�ʐX�щ]<?#J�*� 	�<I2<��J0=�"!�'�2�cg��R�g�7EB��Մ3��H�k�;u(q3U35W�:܋<�2��X����r�$wY��Ϡ�j^�m&����-�AC�����(io	�crU�k�Kޡ�(q2�������zU�H/�3�#�g��7��AB�7�!\4gJ�	 �4�ܟ@NW�o�_.O=��p.��y�7�6	��� �)�
�����Y�a�ӣ�l�g��
�+k�mU�#՘o�8SE��J�P��__?��TM���4��'hZx���&:lk����*5�1b=��T?�{���v�%Iä3��m6֫~�U�&Ɠr0ز]`��G�0��%�#�mw��=3���Q�c��R�T2�~���D����~S8�~j�7���l$��=4 ��2"��[aS�H���J�J9���wt.f���1���v2~����c�GUw��j�[C����Zj�R�y�?$%�b����-���[�ui�M��q?v�
B�1��)�"�^�i���/�d.~�������} T��`��|%�n�n6���9� D���b� �S��N>$�a�Ek�&}�R���b����d|�H�=�D���
�H%��5�Z����ǇQ@I�xp-n��r��η�)P�t���7����˵��h��|"� �|���@�n���E�-��L��"{�FS�Fe����}CP1�;��ꤶ]Kki���b����:�5G鷹��3�����HǮ���}� ���ӊ�o��\A ,����`����TUcH��J�A� ��D�Y�7�*�"No��ɾKRE�0�Ȳ�у*�Rtr�4{�W��4呱 \?fq��q&�������}bb[R���I'~N,t?J��,Zt�G5,	���`�b�i�t�2O��̀r.d���a���[�Zc2\􊜘)��'��#(�<�#��V�S�2�<B'��]O"XZC���G����4_c/�KU]�	*���k�~�`I*�bB8�Kiz_˯ㆺ���;*�K�<�N��pm_ �A�H�RoiOb�$8븵i�l�D� ��eR��W�[
��5&���g��i����u#[��H\�j�:��oU
�%oQ�(i�2�:h+��ل�Oc�U������$� �����)���K4�q|B�ْ��4�����Zx�t`��o�j
�]�9+�G��EJ��R��[߭)���*���LߒJ��t��������_5�V���j���g��K�Xu�q�UQm�#�)�S�$���� �%pN�L��C���&��S3ۀj;��������������J�}�CH7���Cy�}���	 R�S�%�â5q�uc�퍸��+�z9���,W7@Ɲ-�a%�$E�?�_7O>u�ޮ�#��[�W�2)��
�8��=ù>��/�A�tY柺�v75q��^�<x ���