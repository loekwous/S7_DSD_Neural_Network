��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�xW[$�t �T(ڼ�J����(��)BkU���ˢ��2	 ��neG��^=���@���V�ؓt3tk�+��Xه�_(��J���"z��ݗ�#��_®Up\��o�gC���'}�W��4�f׈@��uH�;�`w��3u�s5�A�J�R`��kٶ�B}ʍ~Z��SCT��ᎡUz�s�ȇ5�&�֚�^���o+�++���� @�nB\ie���`Z�5Uw�2@T�x��gA��\U��d
:t�����p�w�s�C�SP�ۥ���͈KP�m���f��3rXj0�� c�7C0C�AԢ���m��Eʨ_�����R��;�. ����թ�ύ�%5�-�F�fWZ�c~��_"�d�0�]L�����8;�(�O�Oq�=v�Iz�H����k��c��nv�њy�S����rDh8x7�J��[2G����-�#{�11�iS�V�VV��	��;[��ag�[icjՖ��Q=��ѱ�~�pd�H��|oU洞�(�D�=�.�5lXAf����R�A�
1�(�>wERIAK@�-���0�â��A�(�i���IJ�c$�����OĢc�Ui;�,`y^mj��W��6�����8#�qg�D�?����]���_�s�L�Ɩ/&{+�n$bVjV����.N��W��hGҭ�lL�?��ر#s���A�Ml�#纠W/v��QB5s!�gd��u ��[.�[L���,�+{f~�"�Ư���?�v��U�4�O,�����a/2����F�V�6�H��*���B����\ \�+��5(���<�0�G\b��V3)�����ҙ�y���]�k�t���=� e6W�8@ӥ�[�]"�>n�bW�/���Г\��z
�T��&����	���t�^�|hwRϳ(5:�{P~_�y�P`��r��v�S�yIn�;� �Vq��K>����&��ib5����Ѥ,&]}<ץ}�H�^{�Ž�V�f�S���A�DP�l�#��dB1鰌�z���V�6������Nޞ[������	�%� ~'i��i��Ә��7k���a��u�����,@V�� ՆgB��o��/���$�l��$�Οh�]3eOp�*���T��ij��-�b�cN�
2�6ۦ[�e�.�|�k�k/u9ޫ�X�����u��W����JP��r=Do{��³Y~�U>Zͣ ���Sa��l��w�-�0�L�O�G�H�h\���&6�{��W=:�K2h�f�LFD&��ϥ1���d->H�9��j,E���b���]�D���!�o@QS�80��O���F�(����j�\N�[X���7�L"�!y��\l�ɳh!�I��6?���"��5�G��TS�^גg��i��7rO����| �b�=|.Jx�O$�.�-Vh7����d�<Z�����s�5EQ�&�{?ey]"Ϛ��!����).W��vW+�C*�2[��_�Բ��,�Ed�� rZ�I��M�΁�?e0�)�ݻ�!�-o� ����?Y�̕Z�=�s���[I&��H-�s
\�3Fb?��q{�������ź=SnI�7jl~���I%0m�	���FācK�FF�!SA�`�rfA��C���@_fYv��sh3
��.�� JXF�~�%Ô{?��u�W\�i�b2�V�����]�4�-!����`�Q:�sI�Z�)��t~+��!8�8Κ�TB��tU���=�����2%�lhx8N���
y=Ğ�<�.:�	F���J�N�����Uq��bو��E�%�aw��,��2\X��sa��/[Oҧ��7z�S�{���P�7�N��R|]��|��E�������K�̦ZK� �݁��D�	�8@����NU��ޘJ$f�g|uD�Lb��&��b�������=�e9_��W��Qg���%��M�BQg[��I�dR�"+d�,Ҩ�Xś+������44}-9.��W�������8��vk��{�7�����eKn�������g��Ydu��ڲ+�l!�Ը�`�X��9�^�{G1��鴶U[����KѸ��Z�9�����!'���-_q��zȑ��d��)'�=�h�8_B����;�!�����R4��}A^5��c�kyeö�c��2 VO�������0��,%�*����Ю������Q8�%ۨr��U@���d���W��Vq�al��`B�ె�ԣ��m��	�*������p�����9�J�U�+qZ֯�C�W<��HA��"4y�(}��
z!��yQ�@���܀g�M�Z���A�'Dy�����O�d*�%/���$8Y�2:t}�qj嬏nR�����	��%�����Ư��A�K|�qd���P\�t��(`���?t�4�*o��D���"m�{C�I��7�~�\t0�ԅU���Q�]m��$JB[iPm@uhO��Rf�\u�)n��)��n����b��J��!]��k�z�Th���h�E��X�(`�5�x���z�d�`�S�䪷����|`��ꟃPɎWQ�e0���0j�=lWJ��7bޱ��k?&�͜cڳ=�w}�7�g�U�����[ˉ�*��=�$I�̊Ԑ#b���Q)X�Q��x)D('���8�8Q0���H�YYֽ,�?�}�Q���q/F"�k�)MEu�8O�o���KC�,� X��$ZTЯ�p���T� �6�!P��V)@Ǣ%��� ]���(&�Kp��q|�cc$E.�}8�gK��R*�������߈��Ί��Iܟi��t3%�l�v�"�6�F����]�0�j�����Kf�CD˾`���A\�g�9	&4Ӈ�^��%sm��_i	�.�!d��ꉸndS&�^k,6:%y��Q3<7� t����0ѫ�����?���?������B
�V1P���+(v��,ۖ�9D2�\�'T�h�&g��޵���8�	^����ݭ�W?��{���9f oI=Z?8qy��п�깫i�*˚\��̿T��OS6r �a��~���U�Aѻ�I�"�6f�/~������Y����7;!����`@�)�����T�d�ݽ�i?ץ9b��ݝD]s���J��A�%5b����Ҙ_Nf&���缐�Fb�����!oQ�]B]u����L�4�Э�>Qq}��$��	a�<w��=�ܵLo��3��dna��8UR�_,r��o��G��[��,_X���_��s���J��d��ͽ�?\��O��@QK�@�.����GoDΗ%=Ix�Q���1l\��c��>�1��/q���p�ɺ�ll��洲l��]��\�~Ԥ8R�l�=�Pc��.".Ҝ�T�G�=�T\0 g��V	E0\�$��x1�¾�7[,�|�u�$
F��P���Z9[�ŧ#�C
5�4<Z�C�x���AV��9��
�n�MЊ�l�1�T��kpڪ�{B��On��&�5���%j�d@���B��d�2���%˴�̃�g�^��K*�=�XM��Uħ�_���+�T�6��=���^C��e�o;�����`�2D�I��ğe�)�,D�mZ]�NP�3FА!3�K�֘�M,u��AT�~�E)�Ȕ;;Ho�1�+��*��4���邝��C��Lm�@l1_��q���g�k��خ����o_�Kr8��qbw�v�1[t4��UJ��<�wSr�};�H�"_®�'����5<��9��Cs/q��f�y,�b�Y�O`#�g������h`�hH&��_T�_�v��������,R��M��`�Y ��'�r������S�tUԷ��+T����X,)�U~< �/Qu�h���`�!<1���78�ͪ�����9���]���&t�Pa**�#�mx4����p�������43�N��Cl���x��*����,�{'�O~�_�01�����|e��z���Ю+��1�	��a�Y�VZ�܋0���h��.�-��X�5�m�W�d���TRُ�e
\��
��{�^=V5+'�$�"]wۂѻP=JC��;�b`?ڔ
���m�� <�^;���q*;e��� F�/�<��=&
S��;�p��g��!�2��nYʴ)�a����Q���ݫ[��r�8�dS�jQXSĥA�K�`�R�"D�����j@yǒEkL����)�U8��sm�#Z���?��<&�m�#��,u�.���"&2?eR^�[�&�nECct9��S�	C�>Ѓ��f�2A�Z����7`��$��K�
5��|o ��s�PZYSb0wsNSp͌i.��>1��sZ{���c��YC����Q�O� T�ﶈ+{{J�؀���v-(�Qߋs�xe���Rm�Pp�!�,8u������m"����"�z�@�߈��Һ�D9&o�~����u���#��pg��C�V��)���l'��{���.��Y
�T�/Z�f΍V���!�.�@�fCi�T����5�V���f����C�,���- ���A�֟��(��R��ooլJ���Kge_�Eq5~�M�8X�\�!�{�+ʛ �k8Ը�J�l66������x]����=E�󀞊ꧾ�<���O����"m ����NP��j1"-U�a��Y��yt���0����o�ceW��Uw�ߺeW��{�����YSڧ�4�#��X���+>o�7KB&����Kz'�W
� N�n�k�΃�.-6����Y0�Ɛ?g�JN�_X[��$�9�g񦃐��^�3:$n��g	�Rssj�s7w-BDs��-"�\%�S�N�_���j��i��ֱ�/�ً6�Ʒ*��K�qĭ�ų(��9��.����M?{=��ws\k�,;�t�V]�n�\�D�U�.CEJ��I���X���R�$ҧ���&�$?FD��߶���~�]��jhERxLȶy�'.oZ���[),i��,�3U�X�y�:^x;侢T[$��l�C��k����d��%}����;6�GbJ�4`�1��g��QR?�c`�1
������ֵ�l��,�|>n��Q��d��6v<��/���4���s��L�ʲ���%���&�y�k�h0~����%�\3�u�qG�?B���.'�1���4�5<����a����8B��Hׁ���"͑�0ç%�2���!6q����rq�	�G��l| $:�ή}��%�C��'4��Z.�aQ_] ���%����W]��q���m�Np�rK����]��k�k �V��*lB��ϙMm�_Lf�����C�qO�?A��+>~~]�j�ȇs����q�z�Y~�~{��N����ʼ~��ciЪHxJ2�~j�=<�{�hM`���qc���e6	o�������lot)j����ɟ�\T/���X;a�